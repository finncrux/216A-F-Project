module Image_Classifier ( 
 input clk, 
 input GlobalReset, 
 input Input_Valid,
 input [18:0] Wgt_0_0, // sfix19_En18 
  input [18:0] Wgt_0_1, // sfix19_En18 
  input [18:0] Wgt_0_2, // sfix19_En18 
  input [18:0] Wgt_0_3, // sfix19_En18 
  input [18:0] Wgt_0_4, // sfix19_En18 
  input [18:0] Wgt_0_5, // sfix19_En18 
  input [18:0] Wgt_0_6, // sfix19_En18 
  input [18:0] Wgt_0_7, // sfix19_En18 
  input [18:0] Wgt_0_8, // sfix19_En18 
  input [18:0] Wgt_0_9, // sfix19_En18 
  input [18:0] Wgt_0_10, // sfix19_En18 
  input [18:0] Wgt_0_11, // sfix19_En18 
  input [18:0] Wgt_0_12, // sfix19_En18 
  input [18:0] Wgt_0_13, // sfix19_En18 
  input [18:0] Wgt_0_14, // sfix19_En18 
  input [18:0] Wgt_0_15, // sfix19_En18 
  input [18:0] Wgt_0_16, // sfix19_En18 
  input [18:0] Wgt_0_17, // sfix19_En18 
  input [18:0] Wgt_0_18, // sfix19_En18 
  input [18:0] Wgt_0_19, // sfix19_En18 
  input [18:0] Wgt_0_20, // sfix19_En18 
  input [18:0] Wgt_0_21, // sfix19_En18 
  input [18:0] Wgt_0_22, // sfix19_En18 
  input [18:0] Wgt_0_23, // sfix19_En18 
  input [18:0] Wgt_0_24, // sfix19_En18 
  input [18:0] Wgt_0_25, // sfix19_En18 
  input [18:0] Wgt_0_26, // sfix19_En18 
  input [18:0] Wgt_0_27, // sfix19_En18 
  input [18:0] Wgt_0_28, // sfix19_En18 
  input [18:0] Wgt_0_29, // sfix19_En18 
  input [18:0] Wgt_0_30, // sfix19_En18 
  input [18:0] Wgt_0_31, // sfix19_En18 
  input [18:0] Wgt_0_32, // sfix19_En18 
  input [18:0] Wgt_0_33, // sfix19_En18 
  input [18:0] Wgt_0_34, // sfix19_En18 
  input [18:0] Wgt_0_35, // sfix19_En18 
  input [18:0] Wgt_0_36, // sfix19_En18 
  input [18:0] Wgt_0_37, // sfix19_En18 
  input [18:0] Wgt_0_38, // sfix19_En18 
  input [18:0] Wgt_0_39, // sfix19_En18 
  input [18:0] Wgt_0_40, // sfix19_En18 
  input [18:0] Wgt_0_41, // sfix19_En18 
  input [18:0] Wgt_0_42, // sfix19_En18 
  input [18:0] Wgt_0_43, // sfix19_En18 
  input [18:0] Wgt_0_44, // sfix19_En18 
  input [18:0] Wgt_0_45, // sfix19_En18 
  input [18:0] Wgt_0_46, // sfix19_En18 
  input [18:0] Wgt_0_47, // sfix19_En18 
  input [18:0] Wgt_0_48, // sfix19_En18 
  input [18:0] Wgt_0_49, // sfix19_En18 
  input [18:0] Wgt_0_50, // sfix19_En18 
  input [18:0] Wgt_0_51, // sfix19_En18 
  input [18:0] Wgt_0_52, // sfix19_En18 
  input [18:0] Wgt_0_53, // sfix19_En18 
  input [18:0] Wgt_0_54, // sfix19_En18 
  input [18:0] Wgt_0_55, // sfix19_En18 
  input [18:0] Wgt_0_56, // sfix19_En18 
  input [18:0] Wgt_0_57, // sfix19_En18 
  input [18:0] Wgt_0_58, // sfix19_En18 
  input [18:0] Wgt_0_59, // sfix19_En18 
  input [18:0] Wgt_0_60, // sfix19_En18 
  input [18:0] Wgt_0_61, // sfix19_En18 
  input [18:0] Wgt_0_62, // sfix19_En18 
  input [18:0] Wgt_0_63, // sfix19_En18 
  input [18:0] Wgt_0_64, // sfix19_En18 
  input [18:0] Wgt_0_65, // sfix19_En18 
  input [18:0] Wgt_0_66, // sfix19_En18 
  input [18:0] Wgt_0_67, // sfix19_En18 
  input [18:0] Wgt_0_68, // sfix19_En18 
  input [18:0] Wgt_0_69, // sfix19_En18 
  input [18:0] Wgt_0_70, // sfix19_En18 
  input [18:0] Wgt_0_71, // sfix19_En18 
  input [18:0] Wgt_0_72, // sfix19_En18 
  input [18:0] Wgt_0_73, // sfix19_En18 
  input [18:0] Wgt_0_74, // sfix19_En18 
  input [18:0] Wgt_0_75, // sfix19_En18 
  input [18:0] Wgt_0_76, // sfix19_En18 
  input [18:0] Wgt_0_77, // sfix19_En18 
  input [18:0] Wgt_0_78, // sfix19_En18 
  input [18:0] Wgt_0_79, // sfix19_En18 
  input [18:0] Wgt_0_80, // sfix19_En18 
  input [18:0] Wgt_0_81, // sfix19_En18 
  input [18:0] Wgt_0_82, // sfix19_En18 
  input [18:0] Wgt_0_83, // sfix19_En18 
  input [18:0] Wgt_0_84, // sfix19_En18 
  input [18:0] Wgt_0_85, // sfix19_En18 
  input [18:0] Wgt_0_86, // sfix19_En18 
  input [18:0] Wgt_0_87, // sfix19_En18 
  input [18:0] Wgt_0_88, // sfix19_En18 
  input [18:0] Wgt_0_89, // sfix19_En18 
  input [18:0] Wgt_0_90, // sfix19_En18 
  input [18:0] Wgt_0_91, // sfix19_En18 
  input [18:0] Wgt_0_92, // sfix19_En18 
  input [18:0] Wgt_0_93, // sfix19_En18 
  input [18:0] Wgt_0_94, // sfix19_En18 
  input [18:0] Wgt_0_95, // sfix19_En18 
  input [18:0] Wgt_0_96, // sfix19_En18 
  input [18:0] Wgt_0_97, // sfix19_En18 
  input [18:0] Wgt_0_98, // sfix19_En18 
  input [18:0] Wgt_0_99, // sfix19_En18 
  input [18:0] Wgt_0_100, // sfix19_En18 
  input [18:0] Wgt_0_101, // sfix19_En18 
  input [18:0] Wgt_0_102, // sfix19_En18 
  input [18:0] Wgt_0_103, // sfix19_En18 
  input [18:0] Wgt_0_104, // sfix19_En18 
  input [18:0] Wgt_0_105, // sfix19_En18 
  input [18:0] Wgt_0_106, // sfix19_En18 
  input [18:0] Wgt_0_107, // sfix19_En18 
  input [18:0] Wgt_0_108, // sfix19_En18 
  input [18:0] Wgt_0_109, // sfix19_En18 
  input [18:0] Wgt_0_110, // sfix19_En18 
  input [18:0] Wgt_0_111, // sfix19_En18 
  input [18:0] Wgt_0_112, // sfix19_En18 
  input [18:0] Wgt_0_113, // sfix19_En18 
  input [18:0] Wgt_0_114, // sfix19_En18 
  input [18:0] Wgt_0_115, // sfix19_En18 
  input [18:0] Wgt_0_116, // sfix19_En18 
  input [18:0] Wgt_0_117, // sfix19_En18 
  input [18:0] Wgt_0_118, // sfix19_En18 
  input [18:0] Wgt_0_119, // sfix19_En18 
  input [18:0] Wgt_0_120, // sfix19_En18 
  input [18:0] Wgt_0_121, // sfix19_En18 
  input [18:0] Wgt_0_122, // sfix19_En18 
  input [18:0] Wgt_0_123, // sfix19_En18 
  input [18:0] Wgt_0_124, // sfix19_En18 
  input [18:0] Wgt_0_125, // sfix19_En18 
  input [18:0] Wgt_0_126, // sfix19_En18 
  input [18:0] Wgt_0_127, // sfix19_En18 
  input [18:0] Wgt_0_128, // sfix19_En18 
  input [18:0] Wgt_0_129, // sfix19_En18 
  input [18:0] Wgt_0_130, // sfix19_En18 
  input [18:0] Wgt_0_131, // sfix19_En18 
  input [18:0] Wgt_0_132, // sfix19_En18 
  input [18:0] Wgt_0_133, // sfix19_En18 
  input [18:0] Wgt_0_134, // sfix19_En18 
  input [18:0] Wgt_0_135, // sfix19_En18 
  input [18:0] Wgt_0_136, // sfix19_En18 
  input [18:0] Wgt_0_137, // sfix19_En18 
  input [18:0] Wgt_0_138, // sfix19_En18 
  input [18:0] Wgt_0_139, // sfix19_En18 
  input [18:0] Wgt_0_140, // sfix19_En18 
  input [18:0] Wgt_0_141, // sfix19_En18 
  input [18:0] Wgt_0_142, // sfix19_En18 
  input [18:0] Wgt_0_143, // sfix19_En18 
  input [18:0] Wgt_0_144, // sfix19_En18 
  input [18:0] Wgt_0_145, // sfix19_En18 
  input [18:0] Wgt_0_146, // sfix19_En18 
  input [18:0] Wgt_0_147, // sfix19_En18 
  input [18:0] Wgt_0_148, // sfix19_En18 
  input [18:0] Wgt_0_149, // sfix19_En18 
  input [18:0] Wgt_0_150, // sfix19_En18 
  input [18:0] Wgt_0_151, // sfix19_En18 
  input [18:0] Wgt_0_152, // sfix19_En18 
  input [18:0] Wgt_0_153, // sfix19_En18 
  input [18:0] Wgt_0_154, // sfix19_En18 
  input [18:0] Wgt_0_155, // sfix19_En18 
  input [18:0] Wgt_0_156, // sfix19_En18 
  input [18:0] Wgt_0_157, // sfix19_En18 
  input [18:0] Wgt_0_158, // sfix19_En18 
  input [18:0] Wgt_0_159, // sfix19_En18 
  input [18:0] Wgt_0_160, // sfix19_En18 
  input [18:0] Wgt_0_161, // sfix19_En18 
  input [18:0] Wgt_0_162, // sfix19_En18 
  input [18:0] Wgt_0_163, // sfix19_En18 
  input [18:0] Wgt_0_164, // sfix19_En18 
  input [18:0] Wgt_0_165, // sfix19_En18 
  input [18:0] Wgt_0_166, // sfix19_En18 
  input [18:0] Wgt_0_167, // sfix19_En18 
  input [18:0] Wgt_0_168, // sfix19_En18 
  input [18:0] Wgt_0_169, // sfix19_En18 
  input [18:0] Wgt_0_170, // sfix19_En18 
  input [18:0] Wgt_0_171, // sfix19_En18 
  input [18:0] Wgt_0_172, // sfix19_En18 
  input [18:0] Wgt_0_173, // sfix19_En18 
  input [18:0] Wgt_0_174, // sfix19_En18 
  input [18:0] Wgt_0_175, // sfix19_En18 
  input [18:0] Wgt_0_176, // sfix19_En18 
  input [18:0] Wgt_0_177, // sfix19_En18 
  input [18:0] Wgt_0_178, // sfix19_En18 
  input [18:0] Wgt_0_179, // sfix19_En18 
  input [18:0] Wgt_0_180, // sfix19_En18 
  input [18:0] Wgt_0_181, // sfix19_En18 
  input [18:0] Wgt_0_182, // sfix19_En18 
  input [18:0] Wgt_0_183, // sfix19_En18 
  input [18:0] Wgt_0_184, // sfix19_En18 
  input [18:0] Wgt_0_185, // sfix19_En18 
  input [18:0] Wgt_0_186, // sfix19_En18 
  input [18:0] Wgt_0_187, // sfix19_En18 
  input [18:0] Wgt_0_188, // sfix19_En18 
  input [18:0] Wgt_0_189, // sfix19_En18 
  input [18:0] Wgt_0_190, // sfix19_En18 
  input [18:0] Wgt_0_191, // sfix19_En18 
  input [18:0] Wgt_0_192, // sfix19_En18 
  input [18:0] Wgt_0_193, // sfix19_En18 
  input [18:0] Wgt_0_194, // sfix19_En18 
  input [18:0] Wgt_0_195, // sfix19_En18 
  input [18:0] Wgt_0_196, // sfix19_En18 
  input [18:0] Wgt_0_197, // sfix19_En18 
  input [18:0] Wgt_0_198, // sfix19_En18 
  input [18:0] Wgt_0_199, // sfix19_En18 
  input [18:0] Wgt_0_200, // sfix19_En18 
  input [18:0] Wgt_0_201, // sfix19_En18 
  input [18:0] Wgt_0_202, // sfix19_En18 
  input [18:0] Wgt_0_203, // sfix19_En18 
  input [18:0] Wgt_0_204, // sfix19_En18 
  input [18:0] Wgt_0_205, // sfix19_En18 
  input [18:0] Wgt_0_206, // sfix19_En18 
  input [18:0] Wgt_0_207, // sfix19_En18 
  input [18:0] Wgt_0_208, // sfix19_En18 
  input [18:0] Wgt_0_209, // sfix19_En18 
  input [18:0] Wgt_0_210, // sfix19_En18 
  input [18:0] Wgt_0_211, // sfix19_En18 
  input [18:0] Wgt_0_212, // sfix19_En18 
  input [18:0] Wgt_0_213, // sfix19_En18 
  input [18:0] Wgt_0_214, // sfix19_En18 
  input [18:0] Wgt_0_215, // sfix19_En18 
  input [18:0] Wgt_0_216, // sfix19_En18 
  input [18:0] Wgt_0_217, // sfix19_En18 
  input [18:0] Wgt_0_218, // sfix19_En18 
  input [18:0] Wgt_0_219, // sfix19_En18 
  input [18:0] Wgt_0_220, // sfix19_En18 
  input [18:0] Wgt_0_221, // sfix19_En18 
  input [18:0] Wgt_0_222, // sfix19_En18 
  input [18:0] Wgt_0_223, // sfix19_En18 
  input [18:0] Wgt_0_224, // sfix19_En18 
  input [18:0] Wgt_0_225, // sfix19_En18 
  input [18:0] Wgt_0_226, // sfix19_En18 
  input [18:0] Wgt_0_227, // sfix19_En18 
  input [18:0] Wgt_0_228, // sfix19_En18 
  input [18:0] Wgt_0_229, // sfix19_En18 
  input [18:0] Wgt_0_230, // sfix19_En18 
  input [18:0] Wgt_0_231, // sfix19_En18 
  input [18:0] Wgt_0_232, // sfix19_En18 
  input [18:0] Wgt_0_233, // sfix19_En18 
  input [18:0] Wgt_0_234, // sfix19_En18 
  input [18:0] Wgt_0_235, // sfix19_En18 
  input [18:0] Wgt_0_236, // sfix19_En18 
  input [18:0] Wgt_0_237, // sfix19_En18 
  input [18:0] Wgt_0_238, // sfix19_En18 
  input [18:0] Wgt_0_239, // sfix19_En18 
  input [18:0] Wgt_0_240, // sfix19_En18 
  input [18:0] Wgt_0_241, // sfix19_En18 
  input [18:0] Wgt_0_242, // sfix19_En18 
  input [18:0] Wgt_0_243, // sfix19_En18 
  input [18:0] Wgt_0_244, // sfix19_En18 
  input [18:0] Wgt_0_245, // sfix19_En18 
  input [18:0] Wgt_0_246, // sfix19_En18 
  input [18:0] Wgt_0_247, // sfix19_En18 
  input [18:0] Wgt_0_248, // sfix19_En18 
  input [18:0] Wgt_0_249, // sfix19_En18 
  input [18:0] Wgt_0_250, // sfix19_En18 
  input [18:0] Wgt_0_251, // sfix19_En18 
  input [18:0] Wgt_0_252, // sfix19_En18 
  input [18:0] Wgt_0_253, // sfix19_En18 
  input [18:0] Wgt_0_254, // sfix19_En18 
  input [18:0] Wgt_0_255, // sfix19_En18 
  input [18:0] Wgt_0_256, // sfix19_En18 
  input [18:0] Wgt_0_257, // sfix19_En18 
  input [18:0] Wgt_0_258, // sfix19_En18 
  input [18:0] Wgt_0_259, // sfix19_En18 
  input [18:0] Wgt_0_260, // sfix19_En18 
  input [18:0] Wgt_0_261, // sfix19_En18 
  input [18:0] Wgt_0_262, // sfix19_En18 
  input [18:0] Wgt_0_263, // sfix19_En18 
  input [18:0] Wgt_0_264, // sfix19_En18 
  input [18:0] Wgt_0_265, // sfix19_En18 
  input [18:0] Wgt_0_266, // sfix19_En18 
  input [18:0] Wgt_0_267, // sfix19_En18 
  input [18:0] Wgt_0_268, // sfix19_En18 
  input [18:0] Wgt_0_269, // sfix19_En18 
  input [18:0] Wgt_0_270, // sfix19_En18 
  input [18:0] Wgt_0_271, // sfix19_En18 
  input [18:0] Wgt_0_272, // sfix19_En18 
  input [18:0] Wgt_0_273, // sfix19_En18 
  input [18:0] Wgt_0_274, // sfix19_En18 
  input [18:0] Wgt_0_275, // sfix19_En18 
  input [18:0] Wgt_0_276, // sfix19_En18 
  input [18:0] Wgt_0_277, // sfix19_En18 
  input [18:0] Wgt_0_278, // sfix19_En18 
  input [18:0] Wgt_0_279, // sfix19_En18 
  input [18:0] Wgt_0_280, // sfix19_En18 
  input [18:0] Wgt_0_281, // sfix19_En18 
  input [18:0] Wgt_0_282, // sfix19_En18 
  input [18:0] Wgt_0_283, // sfix19_En18 
  input [18:0] Wgt_0_284, // sfix19_En18 
  input [18:0] Wgt_0_285, // sfix19_En18 
  input [18:0] Wgt_0_286, // sfix19_En18 
  input [18:0] Wgt_0_287, // sfix19_En18 
  input [18:0] Wgt_0_288, // sfix19_En18 
  input [18:0] Wgt_0_289, // sfix19_En18 
  input [18:0] Wgt_0_290, // sfix19_En18 
  input [18:0] Wgt_0_291, // sfix19_En18 
  input [18:0] Wgt_0_292, // sfix19_En18 
  input [18:0] Wgt_0_293, // sfix19_En18 
  input [18:0] Wgt_0_294, // sfix19_En18 
  input [18:0] Wgt_0_295, // sfix19_En18 
  input [18:0] Wgt_0_296, // sfix19_En18 
  input [18:0] Wgt_0_297, // sfix19_En18 
  input [18:0] Wgt_0_298, // sfix19_En18 
  input [18:0] Wgt_0_299, // sfix19_En18 
  input [18:0] Wgt_0_300, // sfix19_En18 
  input [18:0] Wgt_0_301, // sfix19_En18 
  input [18:0] Wgt_0_302, // sfix19_En18 
  input [18:0] Wgt_0_303, // sfix19_En18 
  input [18:0] Wgt_0_304, // sfix19_En18 
  input [18:0] Wgt_0_305, // sfix19_En18 
  input [18:0] Wgt_0_306, // sfix19_En18 
  input [18:0] Wgt_0_307, // sfix19_En18 
  input [18:0] Wgt_0_308, // sfix19_En18 
  input [18:0] Wgt_0_309, // sfix19_En18 
  input [18:0] Wgt_0_310, // sfix19_En18 
  input [18:0] Wgt_0_311, // sfix19_En18 
  input [18:0] Wgt_0_312, // sfix19_En18 
  input [18:0] Wgt_0_313, // sfix19_En18 
  input [18:0] Wgt_0_314, // sfix19_En18 
  input [18:0] Wgt_0_315, // sfix19_En18 
  input [18:0] Wgt_0_316, // sfix19_En18 
  input [18:0] Wgt_0_317, // sfix19_En18 
  input [18:0] Wgt_0_318, // sfix19_En18 
  input [18:0] Wgt_0_319, // sfix19_En18 
  input [18:0] Wgt_0_320, // sfix19_En18 
  input [18:0] Wgt_0_321, // sfix19_En18 
  input [18:0] Wgt_0_322, // sfix19_En18 
  input [18:0] Wgt_0_323, // sfix19_En18 
  input [18:0] Wgt_0_324, // sfix19_En18 
  input [18:0] Wgt_0_325, // sfix19_En18 
  input [18:0] Wgt_0_326, // sfix19_En18 
  input [18:0] Wgt_0_327, // sfix19_En18 
  input [18:0] Wgt_0_328, // sfix19_En18 
  input [18:0] Wgt_0_329, // sfix19_En18 
  input [18:0] Wgt_0_330, // sfix19_En18 
  input [18:0] Wgt_0_331, // sfix19_En18 
  input [18:0] Wgt_0_332, // sfix19_En18 
  input [18:0] Wgt_0_333, // sfix19_En18 
  input [18:0] Wgt_0_334, // sfix19_En18 
  input [18:0] Wgt_0_335, // sfix19_En18 
  input [18:0] Wgt_0_336, // sfix19_En18 
  input [18:0] Wgt_0_337, // sfix19_En18 
  input [18:0] Wgt_0_338, // sfix19_En18 
  input [18:0] Wgt_0_339, // sfix19_En18 
  input [18:0] Wgt_0_340, // sfix19_En18 
  input [18:0] Wgt_0_341, // sfix19_En18 
  input [18:0] Wgt_0_342, // sfix19_En18 
  input [18:0] Wgt_0_343, // sfix19_En18 
  input [18:0] Wgt_0_344, // sfix19_En18 
  input [18:0] Wgt_0_345, // sfix19_En18 
  input [18:0] Wgt_0_346, // sfix19_En18 
  input [18:0] Wgt_0_347, // sfix19_En18 
  input [18:0] Wgt_0_348, // sfix19_En18 
  input [18:0] Wgt_0_349, // sfix19_En18 
  input [18:0] Wgt_0_350, // sfix19_En18 
  input [18:0] Wgt_0_351, // sfix19_En18 
  input [18:0] Wgt_0_352, // sfix19_En18 
  input [18:0] Wgt_0_353, // sfix19_En18 
  input [18:0] Wgt_0_354, // sfix19_En18 
  input [18:0] Wgt_0_355, // sfix19_En18 
  input [18:0] Wgt_0_356, // sfix19_En18 
  input [18:0] Wgt_0_357, // sfix19_En18 
  input [18:0] Wgt_0_358, // sfix19_En18 
  input [18:0] Wgt_0_359, // sfix19_En18 
  input [18:0] Wgt_0_360, // sfix19_En18 
  input [18:0] Wgt_0_361, // sfix19_En18 
  input [18:0] Wgt_0_362, // sfix19_En18 
  input [18:0] Wgt_0_363, // sfix19_En18 
  input [18:0] Wgt_0_364, // sfix19_En18 
  input [18:0] Wgt_0_365, // sfix19_En18 
  input [18:0] Wgt_0_366, // sfix19_En18 
  input [18:0] Wgt_0_367, // sfix19_En18 
  input [18:0] Wgt_0_368, // sfix19_En18 
  input [18:0] Wgt_0_369, // sfix19_En18 
  input [18:0] Wgt_0_370, // sfix19_En18 
  input [18:0] Wgt_0_371, // sfix19_En18 
  input [18:0] Wgt_0_372, // sfix19_En18 
  input [18:0] Wgt_0_373, // sfix19_En18 
  input [18:0] Wgt_0_374, // sfix19_En18 
  input [18:0] Wgt_0_375, // sfix19_En18 
  input [18:0] Wgt_0_376, // sfix19_En18 
  input [18:0] Wgt_0_377, // sfix19_En18 
  input [18:0] Wgt_0_378, // sfix19_En18 
  input [18:0] Wgt_0_379, // sfix19_En18 
  input [18:0] Wgt_0_380, // sfix19_En18 
  input [18:0] Wgt_0_381, // sfix19_En18 
  input [18:0] Wgt_0_382, // sfix19_En18 
  input [18:0] Wgt_0_383, // sfix19_En18 
  input [18:0] Wgt_0_384, // sfix19_En18 
  input [18:0] Wgt_0_385, // sfix19_En18 
  input [18:0] Wgt_0_386, // sfix19_En18 
  input [18:0] Wgt_0_387, // sfix19_En18 
  input [18:0] Wgt_0_388, // sfix19_En18 
  input [18:0] Wgt_0_389, // sfix19_En18 
  input [18:0] Wgt_0_390, // sfix19_En18 
  input [18:0] Wgt_0_391, // sfix19_En18 
  input [18:0] Wgt_0_392, // sfix19_En18 
  input [18:0] Wgt_0_393, // sfix19_En18 
  input [18:0] Wgt_0_394, // sfix19_En18 
  input [18:0] Wgt_0_395, // sfix19_En18 
  input [18:0] Wgt_0_396, // sfix19_En18 
  input [18:0] Wgt_0_397, // sfix19_En18 
  input [18:0] Wgt_0_398, // sfix19_En18 
  input [18:0] Wgt_0_399, // sfix19_En18 
  input [18:0] Wgt_0_400, // sfix19_En18 
  input [18:0] Wgt_0_401, // sfix19_En18 
  input [18:0] Wgt_0_402, // sfix19_En18 
  input [18:0] Wgt_0_403, // sfix19_En18 
  input [18:0] Wgt_0_404, // sfix19_En18 
  input [18:0] Wgt_0_405, // sfix19_En18 
  input [18:0] Wgt_0_406, // sfix19_En18 
  input [18:0] Wgt_0_407, // sfix19_En18 
  input [18:0] Wgt_0_408, // sfix19_En18 
  input [18:0] Wgt_0_409, // sfix19_En18 
  input [18:0] Wgt_0_410, // sfix19_En18 
  input [18:0] Wgt_0_411, // sfix19_En18 
  input [18:0] Wgt_0_412, // sfix19_En18 
  input [18:0] Wgt_0_413, // sfix19_En18 
  input [18:0] Wgt_0_414, // sfix19_En18 
  input [18:0] Wgt_0_415, // sfix19_En18 
  input [18:0] Wgt_0_416, // sfix19_En18 
  input [18:0] Wgt_0_417, // sfix19_En18 
  input [18:0] Wgt_0_418, // sfix19_En18 
  input [18:0] Wgt_0_419, // sfix19_En18 
  input [18:0] Wgt_0_420, // sfix19_En18 
  input [18:0] Wgt_0_421, // sfix19_En18 
  input [18:0] Wgt_0_422, // sfix19_En18 
  input [18:0] Wgt_0_423, // sfix19_En18 
  input [18:0] Wgt_0_424, // sfix19_En18 
  input [18:0] Wgt_0_425, // sfix19_En18 
  input [18:0] Wgt_0_426, // sfix19_En18 
  input [18:0] Wgt_0_427, // sfix19_En18 
  input [18:0] Wgt_0_428, // sfix19_En18 
  input [18:0] Wgt_0_429, // sfix19_En18 
  input [18:0] Wgt_0_430, // sfix19_En18 
  input [18:0] Wgt_0_431, // sfix19_En18 
  input [18:0] Wgt_0_432, // sfix19_En18 
  input [18:0] Wgt_0_433, // sfix19_En18 
  input [18:0] Wgt_0_434, // sfix19_En18 
  input [18:0] Wgt_0_435, // sfix19_En18 
  input [18:0] Wgt_0_436, // sfix19_En18 
  input [18:0] Wgt_0_437, // sfix19_En18 
  input [18:0] Wgt_0_438, // sfix19_En18 
  input [18:0] Wgt_0_439, // sfix19_En18 
  input [18:0] Wgt_0_440, // sfix19_En18 
  input [18:0] Wgt_0_441, // sfix19_En18 
  input [18:0] Wgt_0_442, // sfix19_En18 
  input [18:0] Wgt_0_443, // sfix19_En18 
  input [18:0] Wgt_0_444, // sfix19_En18 
  input [18:0] Wgt_0_445, // sfix19_En18 
  input [18:0] Wgt_0_446, // sfix19_En18 
  input [18:0] Wgt_0_447, // sfix19_En18 
  input [18:0] Wgt_0_448, // sfix19_En18 
  input [18:0] Wgt_0_449, // sfix19_En18 
  input [18:0] Wgt_0_450, // sfix19_En18 
  input [18:0] Wgt_0_451, // sfix19_En18 
  input [18:0] Wgt_0_452, // sfix19_En18 
  input [18:0] Wgt_0_453, // sfix19_En18 
  input [18:0] Wgt_0_454, // sfix19_En18 
  input [18:0] Wgt_0_455, // sfix19_En18 
  input [18:0] Wgt_0_456, // sfix19_En18 
  input [18:0] Wgt_0_457, // sfix19_En18 
  input [18:0] Wgt_0_458, // sfix19_En18 
  input [18:0] Wgt_0_459, // sfix19_En18 
  input [18:0] Wgt_0_460, // sfix19_En18 
  input [18:0] Wgt_0_461, // sfix19_En18 
  input [18:0] Wgt_0_462, // sfix19_En18 
  input [18:0] Wgt_0_463, // sfix19_En18 
  input [18:0] Wgt_0_464, // sfix19_En18 
  input [18:0] Wgt_0_465, // sfix19_En18 
  input [18:0] Wgt_0_466, // sfix19_En18 
  input [18:0] Wgt_0_467, // sfix19_En18 
  input [18:0] Wgt_0_468, // sfix19_En18 
  input [18:0] Wgt_0_469, // sfix19_En18 
  input [18:0] Wgt_0_470, // sfix19_En18 
  input [18:0] Wgt_0_471, // sfix19_En18 
  input [18:0] Wgt_0_472, // sfix19_En18 
  input [18:0] Wgt_0_473, // sfix19_En18 
  input [18:0] Wgt_0_474, // sfix19_En18 
  input [18:0] Wgt_0_475, // sfix19_En18 
  input [18:0] Wgt_0_476, // sfix19_En18 
  input [18:0] Wgt_0_477, // sfix19_En18 
  input [18:0] Wgt_0_478, // sfix19_En18 
  input [18:0] Wgt_0_479, // sfix19_En18 
  input [18:0] Wgt_0_480, // sfix19_En18 
  input [18:0] Wgt_0_481, // sfix19_En18 
  input [18:0] Wgt_0_482, // sfix19_En18 
  input [18:0] Wgt_0_483, // sfix19_En18 
  input [18:0] Wgt_0_484, // sfix19_En18 
  input [18:0] Wgt_0_485, // sfix19_En18 
  input [18:0] Wgt_0_486, // sfix19_En18 
  input [18:0] Wgt_0_487, // sfix19_En18 
  input [18:0] Wgt_0_488, // sfix19_En18 
  input [18:0] Wgt_0_489, // sfix19_En18 
  input [18:0] Wgt_0_490, // sfix19_En18 
  input [18:0] Wgt_0_491, // sfix19_En18 
  input [18:0] Wgt_0_492, // sfix19_En18 
  input [18:0] Wgt_0_493, // sfix19_En18 
  input [18:0] Wgt_0_494, // sfix19_En18 
  input [18:0] Wgt_0_495, // sfix19_En18 
  input [18:0] Wgt_0_496, // sfix19_En18 
  input [18:0] Wgt_0_497, // sfix19_En18 
  input [18:0] Wgt_0_498, // sfix19_En18 
  input [18:0] Wgt_0_499, // sfix19_En18 
  input [18:0] Wgt_0_500, // sfix19_En18 
  input [18:0] Wgt_0_501, // sfix19_En18 
  input [18:0] Wgt_0_502, // sfix19_En18 
  input [18:0] Wgt_0_503, // sfix19_En18 
  input [18:0] Wgt_0_504, // sfix19_En18 
  input [18:0] Wgt_0_505, // sfix19_En18 
  input [18:0] Wgt_0_506, // sfix19_En18 
  input [18:0] Wgt_0_507, // sfix19_En18 
  input [18:0] Wgt_0_508, // sfix19_En18 
  input [18:0] Wgt_0_509, // sfix19_En18 
  input [18:0] Wgt_0_510, // sfix19_En18 
  input [18:0] Wgt_0_511, // sfix19_En18 
  input [18:0] Wgt_0_512, // sfix19_En18 
  input [18:0] Wgt_0_513, // sfix19_En18 
  input [18:0] Wgt_0_514, // sfix19_En18 
  input [18:0] Wgt_0_515, // sfix19_En18 
  input [18:0] Wgt_0_516, // sfix19_En18 
  input [18:0] Wgt_0_517, // sfix19_En18 
  input [18:0] Wgt_0_518, // sfix19_En18 
  input [18:0] Wgt_0_519, // sfix19_En18 
  input [18:0] Wgt_0_520, // sfix19_En18 
  input [18:0] Wgt_0_521, // sfix19_En18 
  input [18:0] Wgt_0_522, // sfix19_En18 
  input [18:0] Wgt_0_523, // sfix19_En18 
  input [18:0] Wgt_0_524, // sfix19_En18 
  input [18:0] Wgt_0_525, // sfix19_En18 
  input [18:0] Wgt_0_526, // sfix19_En18 
  input [18:0] Wgt_0_527, // sfix19_En18 
  input [18:0] Wgt_0_528, // sfix19_En18 
  input [18:0] Wgt_0_529, // sfix19_En18 
  input [18:0] Wgt_0_530, // sfix19_En18 
  input [18:0] Wgt_0_531, // sfix19_En18 
  input [18:0] Wgt_0_532, // sfix19_En18 
  input [18:0] Wgt_0_533, // sfix19_En18 
  input [18:0] Wgt_0_534, // sfix19_En18 
  input [18:0] Wgt_0_535, // sfix19_En18 
  input [18:0] Wgt_0_536, // sfix19_En18 
  input [18:0] Wgt_0_537, // sfix19_En18 
  input [18:0] Wgt_0_538, // sfix19_En18 
  input [18:0] Wgt_0_539, // sfix19_En18 
  input [18:0] Wgt_0_540, // sfix19_En18 
  input [18:0] Wgt_0_541, // sfix19_En18 
  input [18:0] Wgt_0_542, // sfix19_En18 
  input [18:0] Wgt_0_543, // sfix19_En18 
  input [18:0] Wgt_0_544, // sfix19_En18 
  input [18:0] Wgt_0_545, // sfix19_En18 
  input [18:0] Wgt_0_546, // sfix19_En18 
  input [18:0] Wgt_0_547, // sfix19_En18 
  input [18:0] Wgt_0_548, // sfix19_En18 
  input [18:0] Wgt_0_549, // sfix19_En18 
  input [18:0] Wgt_0_550, // sfix19_En18 
  input [18:0] Wgt_0_551, // sfix19_En18 
  input [18:0] Wgt_0_552, // sfix19_En18 
  input [18:0] Wgt_0_553, // sfix19_En18 
  input [18:0] Wgt_0_554, // sfix19_En18 
  input [18:0] Wgt_0_555, // sfix19_En18 
  input [18:0] Wgt_0_556, // sfix19_En18 
  input [18:0] Wgt_0_557, // sfix19_En18 
  input [18:0] Wgt_0_558, // sfix19_En18 
  input [18:0] Wgt_0_559, // sfix19_En18 
  input [18:0] Wgt_0_560, // sfix19_En18 
  input [18:0] Wgt_0_561, // sfix19_En18 
  input [18:0] Wgt_0_562, // sfix19_En18 
  input [18:0] Wgt_0_563, // sfix19_En18 
  input [18:0] Wgt_0_564, // sfix19_En18 
  input [18:0] Wgt_0_565, // sfix19_En18 
  input [18:0] Wgt_0_566, // sfix19_En18 
  input [18:0] Wgt_0_567, // sfix19_En18 
  input [18:0] Wgt_0_568, // sfix19_En18 
  input [18:0] Wgt_0_569, // sfix19_En18 
  input [18:0] Wgt_0_570, // sfix19_En18 
  input [18:0] Wgt_0_571, // sfix19_En18 
  input [18:0] Wgt_0_572, // sfix19_En18 
  input [18:0] Wgt_0_573, // sfix19_En18 
  input [18:0] Wgt_0_574, // sfix19_En18 
  input [18:0] Wgt_0_575, // sfix19_En18 
  input [18:0] Wgt_0_576, // sfix19_En18 
  input [18:0] Wgt_0_577, // sfix19_En18 
  input [18:0] Wgt_0_578, // sfix19_En18 
  input [18:0] Wgt_0_579, // sfix19_En18 
  input [18:0] Wgt_0_580, // sfix19_En18 
  input [18:0] Wgt_0_581, // sfix19_En18 
  input [18:0] Wgt_0_582, // sfix19_En18 
  input [18:0] Wgt_0_583, // sfix19_En18 
  input [18:0] Wgt_0_584, // sfix19_En18 
  input [18:0] Wgt_0_585, // sfix19_En18 
  input [18:0] Wgt_0_586, // sfix19_En18 
  input [18:0] Wgt_0_587, // sfix19_En18 
  input [18:0] Wgt_0_588, // sfix19_En18 
  input [18:0] Wgt_0_589, // sfix19_En18 
  input [18:0] Wgt_0_590, // sfix19_En18 
  input [18:0] Wgt_0_591, // sfix19_En18 
  input [18:0] Wgt_0_592, // sfix19_En18 
  input [18:0] Wgt_0_593, // sfix19_En18 
  input [18:0] Wgt_0_594, // sfix19_En18 
  input [18:0] Wgt_0_595, // sfix19_En18 
  input [18:0] Wgt_0_596, // sfix19_En18 
  input [18:0] Wgt_0_597, // sfix19_En18 
  input [18:0] Wgt_0_598, // sfix19_En18 
  input [18:0] Wgt_0_599, // sfix19_En18 
  input [18:0] Wgt_0_600, // sfix19_En18 
  input [18:0] Wgt_0_601, // sfix19_En18 
  input [18:0] Wgt_0_602, // sfix19_En18 
  input [18:0] Wgt_0_603, // sfix19_En18 
  input [18:0] Wgt_0_604, // sfix19_En18 
  input [18:0] Wgt_0_605, // sfix19_En18 
  input [18:0] Wgt_0_606, // sfix19_En18 
  input [18:0] Wgt_0_607, // sfix19_En18 
  input [18:0] Wgt_0_608, // sfix19_En18 
  input [18:0] Wgt_0_609, // sfix19_En18 
  input [18:0] Wgt_0_610, // sfix19_En18 
  input [18:0] Wgt_0_611, // sfix19_En18 
  input [18:0] Wgt_0_612, // sfix19_En18 
  input [18:0] Wgt_0_613, // sfix19_En18 
  input [18:0] Wgt_0_614, // sfix19_En18 
  input [18:0] Wgt_0_615, // sfix19_En18 
  input [18:0] Wgt_0_616, // sfix19_En18 
  input [18:0] Wgt_0_617, // sfix19_En18 
  input [18:0] Wgt_0_618, // sfix19_En18 
  input [18:0] Wgt_0_619, // sfix19_En18 
  input [18:0] Wgt_0_620, // sfix19_En18 
  input [18:0] Wgt_0_621, // sfix19_En18 
  input [18:0] Wgt_0_622, // sfix19_En18 
  input [18:0] Wgt_0_623, // sfix19_En18 
  input [18:0] Wgt_0_624, // sfix19_En18 
  input [18:0] Wgt_0_625, // sfix19_En18 
  input [18:0] Wgt_0_626, // sfix19_En18 
  input [18:0] Wgt_0_627, // sfix19_En18 
  input [18:0] Wgt_0_628, // sfix19_En18 
  input [18:0] Wgt_0_629, // sfix19_En18 
  input [18:0] Wgt_0_630, // sfix19_En18 
  input [18:0] Wgt_0_631, // sfix19_En18 
  input [18:0] Wgt_0_632, // sfix19_En18 
  input [18:0] Wgt_0_633, // sfix19_En18 
  input [18:0] Wgt_0_634, // sfix19_En18 
  input [18:0] Wgt_0_635, // sfix19_En18 
  input [18:0] Wgt_0_636, // sfix19_En18 
  input [18:0] Wgt_0_637, // sfix19_En18 
  input [18:0] Wgt_0_638, // sfix19_En18 
  input [18:0] Wgt_0_639, // sfix19_En18 
  input [18:0] Wgt_0_640, // sfix19_En18 
  input [18:0] Wgt_0_641, // sfix19_En18 
  input [18:0] Wgt_0_642, // sfix19_En18 
  input [18:0] Wgt_0_643, // sfix19_En18 
  input [18:0] Wgt_0_644, // sfix19_En18 
  input [18:0] Wgt_0_645, // sfix19_En18 
  input [18:0] Wgt_0_646, // sfix19_En18 
  input [18:0] Wgt_0_647, // sfix19_En18 
  input [18:0] Wgt_0_648, // sfix19_En18 
  input [18:0] Wgt_0_649, // sfix19_En18 
  input [18:0] Wgt_0_650, // sfix19_En18 
  input [18:0] Wgt_0_651, // sfix19_En18 
  input [18:0] Wgt_0_652, // sfix19_En18 
  input [18:0] Wgt_0_653, // sfix19_En18 
  input [18:0] Wgt_0_654, // sfix19_En18 
  input [18:0] Wgt_0_655, // sfix19_En18 
  input [18:0] Wgt_0_656, // sfix19_En18 
  input [18:0] Wgt_0_657, // sfix19_En18 
  input [18:0] Wgt_0_658, // sfix19_En18 
  input [18:0] Wgt_0_659, // sfix19_En18 
  input [18:0] Wgt_0_660, // sfix19_En18 
  input [18:0] Wgt_0_661, // sfix19_En18 
  input [18:0] Wgt_0_662, // sfix19_En18 
  input [18:0] Wgt_0_663, // sfix19_En18 
  input [18:0] Wgt_0_664, // sfix19_En18 
  input [18:0] Wgt_0_665, // sfix19_En18 
  input [18:0] Wgt_0_666, // sfix19_En18 
  input [18:0] Wgt_0_667, // sfix19_En18 
  input [18:0] Wgt_0_668, // sfix19_En18 
  input [18:0] Wgt_0_669, // sfix19_En18 
  input [18:0] Wgt_0_670, // sfix19_En18 
  input [18:0] Wgt_0_671, // sfix19_En18 
  input [18:0] Wgt_0_672, // sfix19_En18 
  input [18:0] Wgt_0_673, // sfix19_En18 
  input [18:0] Wgt_0_674, // sfix19_En18 
  input [18:0] Wgt_0_675, // sfix19_En18 
  input [18:0] Wgt_0_676, // sfix19_En18 
  input [18:0] Wgt_0_677, // sfix19_En18 
  input [18:0] Wgt_0_678, // sfix19_En18 
  input [18:0] Wgt_0_679, // sfix19_En18 
  input [18:0] Wgt_0_680, // sfix19_En18 
  input [18:0] Wgt_0_681, // sfix19_En18 
  input [18:0] Wgt_0_682, // sfix19_En18 
  input [18:0] Wgt_0_683, // sfix19_En18 
  input [18:0] Wgt_0_684, // sfix19_En18 
  input [18:0] Wgt_0_685, // sfix19_En18 
  input [18:0] Wgt_0_686, // sfix19_En18 
  input [18:0] Wgt_0_687, // sfix19_En18 
  input [18:0] Wgt_0_688, // sfix19_En18 
  input [18:0] Wgt_0_689, // sfix19_En18 
  input [18:0] Wgt_0_690, // sfix19_En18 
  input [18:0] Wgt_0_691, // sfix19_En18 
  input [18:0] Wgt_0_692, // sfix19_En18 
  input [18:0] Wgt_0_693, // sfix19_En18 
  input [18:0] Wgt_0_694, // sfix19_En18 
  input [18:0] Wgt_0_695, // sfix19_En18 
  input [18:0] Wgt_0_696, // sfix19_En18 
  input [18:0] Wgt_0_697, // sfix19_En18 
  input [18:0] Wgt_0_698, // sfix19_En18 
  input [18:0] Wgt_0_699, // sfix19_En18 
  input [18:0] Wgt_0_700, // sfix19_En18 
  input [18:0] Wgt_0_701, // sfix19_En18 
  input [18:0] Wgt_0_702, // sfix19_En18 
  input [18:0] Wgt_0_703, // sfix19_En18 
  input [18:0] Wgt_0_704, // sfix19_En18 
  input [18:0] Wgt_0_705, // sfix19_En18 
  input [18:0] Wgt_0_706, // sfix19_En18 
  input [18:0] Wgt_0_707, // sfix19_En18 
  input [18:0] Wgt_0_708, // sfix19_En18 
  input [18:0] Wgt_0_709, // sfix19_En18 
  input [18:0] Wgt_0_710, // sfix19_En18 
  input [18:0] Wgt_0_711, // sfix19_En18 
  input [18:0] Wgt_0_712, // sfix19_En18 
  input [18:0] Wgt_0_713, // sfix19_En18 
  input [18:0] Wgt_0_714, // sfix19_En18 
  input [18:0] Wgt_0_715, // sfix19_En18 
  input [18:0] Wgt_0_716, // sfix19_En18 
  input [18:0] Wgt_0_717, // sfix19_En18 
  input [18:0] Wgt_0_718, // sfix19_En18 
  input [18:0] Wgt_0_719, // sfix19_En18 
  input [18:0] Wgt_0_720, // sfix19_En18 
  input [18:0] Wgt_0_721, // sfix19_En18 
  input [18:0] Wgt_0_722, // sfix19_En18 
  input [18:0] Wgt_0_723, // sfix19_En18 
  input [18:0] Wgt_0_724, // sfix19_En18 
  input [18:0] Wgt_0_725, // sfix19_En18 
  input [18:0] Wgt_0_726, // sfix19_En18 
  input [18:0] Wgt_0_727, // sfix19_En18 
  input [18:0] Wgt_0_728, // sfix19_En18 
  input [18:0] Wgt_0_729, // sfix19_En18 
  input [18:0] Wgt_0_730, // sfix19_En18 
  input [18:0] Wgt_0_731, // sfix19_En18 
  input [18:0] Wgt_0_732, // sfix19_En18 
  input [18:0] Wgt_0_733, // sfix19_En18 
  input [18:0] Wgt_0_734, // sfix19_En18 
  input [18:0] Wgt_0_735, // sfix19_En18 
  input [18:0] Wgt_0_736, // sfix19_En18 
  input [18:0] Wgt_0_737, // sfix19_En18 
  input [18:0] Wgt_0_738, // sfix19_En18 
  input [18:0] Wgt_0_739, // sfix19_En18 
  input [18:0] Wgt_0_740, // sfix19_En18 
  input [18:0] Wgt_0_741, // sfix19_En18 
  input [18:0] Wgt_0_742, // sfix19_En18 
  input [18:0] Wgt_0_743, // sfix19_En18 
  input [18:0] Wgt_0_744, // sfix19_En18 
  input [18:0] Wgt_0_745, // sfix19_En18 
  input [18:0] Wgt_0_746, // sfix19_En18 
  input [18:0] Wgt_0_747, // sfix19_En18 
  input [18:0] Wgt_0_748, // sfix19_En18 
  input [18:0] Wgt_0_749, // sfix19_En18 
  input [18:0] Wgt_0_750, // sfix19_En18 
  input [18:0] Wgt_0_751, // sfix19_En18 
  input [18:0] Wgt_0_752, // sfix19_En18 
  input [18:0] Wgt_0_753, // sfix19_En18 
  input [18:0] Wgt_0_754, // sfix19_En18 
  input [18:0] Wgt_0_755, // sfix19_En18 
  input [18:0] Wgt_0_756, // sfix19_En18 
  input [18:0] Wgt_0_757, // sfix19_En18 
  input [18:0] Wgt_0_758, // sfix19_En18 
  input [18:0] Wgt_0_759, // sfix19_En18 
  input [18:0] Wgt_0_760, // sfix19_En18 
  input [18:0] Wgt_0_761, // sfix19_En18 
  input [18:0] Wgt_0_762, // sfix19_En18 
  input [18:0] Wgt_0_763, // sfix19_En18 
  input [18:0] Wgt_0_764, // sfix19_En18 
  input [18:0] Wgt_0_765, // sfix19_En18 
  input [18:0] Wgt_0_766, // sfix19_En18 
  input [18:0] Wgt_0_767, // sfix19_En18 
  input [18:0] Wgt_0_768, // sfix19_En18 
  input [18:0] Wgt_0_769, // sfix19_En18 
  input [18:0] Wgt_0_770, // sfix19_En18 
  input [18:0] Wgt_0_771, // sfix19_En18 
  input [18:0] Wgt_0_772, // sfix19_En18 
  input [18:0] Wgt_0_773, // sfix19_En18 
  input [18:0] Wgt_0_774, // sfix19_En18 
  input [18:0] Wgt_0_775, // sfix19_En18 
  input [18:0] Wgt_0_776, // sfix19_En18 
  input [18:0] Wgt_0_777, // sfix19_En18 
  input [18:0] Wgt_0_778, // sfix19_En18 
  input [18:0] Wgt_0_779, // sfix19_En18 
  input [18:0] Wgt_0_780, // sfix19_En18 
  input [18:0] Wgt_0_781, // sfix19_En18 
  input [18:0] Wgt_0_782, // sfix19_En18 
  input [18:0] Wgt_0_783, // sfix19_En18 
  input [18:0] Wgt_0_784, // sfix19_En18 
  input [18:0] Wgt_1_0, // sfix19_En18 
  input [18:0] Wgt_1_1, // sfix19_En18 
  input [18:0] Wgt_1_2, // sfix19_En18 
  input [18:0] Wgt_1_3, // sfix19_En18 
  input [18:0] Wgt_1_4, // sfix19_En18 
  input [18:0] Wgt_1_5, // sfix19_En18 
  input [18:0] Wgt_1_6, // sfix19_En18 
  input [18:0] Wgt_1_7, // sfix19_En18 
  input [18:0] Wgt_1_8, // sfix19_En18 
  input [18:0] Wgt_1_9, // sfix19_En18 
  input [18:0] Wgt_1_10, // sfix19_En18 
  input [18:0] Wgt_1_11, // sfix19_En18 
  input [18:0] Wgt_1_12, // sfix19_En18 
  input [18:0] Wgt_1_13, // sfix19_En18 
  input [18:0] Wgt_1_14, // sfix19_En18 
  input [18:0] Wgt_1_15, // sfix19_En18 
  input [18:0] Wgt_1_16, // sfix19_En18 
  input [18:0] Wgt_1_17, // sfix19_En18 
  input [18:0] Wgt_1_18, // sfix19_En18 
  input [18:0] Wgt_1_19, // sfix19_En18 
  input [18:0] Wgt_1_20, // sfix19_En18 
  input [18:0] Wgt_1_21, // sfix19_En18 
  input [18:0] Wgt_1_22, // sfix19_En18 
  input [18:0] Wgt_1_23, // sfix19_En18 
  input [18:0] Wgt_1_24, // sfix19_En18 
  input [18:0] Wgt_1_25, // sfix19_En18 
  input [18:0] Wgt_1_26, // sfix19_En18 
  input [18:0] Wgt_1_27, // sfix19_En18 
  input [18:0] Wgt_1_28, // sfix19_En18 
  input [18:0] Wgt_1_29, // sfix19_En18 
  input [18:0] Wgt_1_30, // sfix19_En18 
  input [18:0] Wgt_1_31, // sfix19_En18 
  input [18:0] Wgt_1_32, // sfix19_En18 
  input [18:0] Wgt_1_33, // sfix19_En18 
  input [18:0] Wgt_1_34, // sfix19_En18 
  input [18:0] Wgt_1_35, // sfix19_En18 
  input [18:0] Wgt_1_36, // sfix19_En18 
  input [18:0] Wgt_1_37, // sfix19_En18 
  input [18:0] Wgt_1_38, // sfix19_En18 
  input [18:0] Wgt_1_39, // sfix19_En18 
  input [18:0] Wgt_1_40, // sfix19_En18 
  input [18:0] Wgt_1_41, // sfix19_En18 
  input [18:0] Wgt_1_42, // sfix19_En18 
  input [18:0] Wgt_1_43, // sfix19_En18 
  input [18:0] Wgt_1_44, // sfix19_En18 
  input [18:0] Wgt_1_45, // sfix19_En18 
  input [18:0] Wgt_1_46, // sfix19_En18 
  input [18:0] Wgt_1_47, // sfix19_En18 
  input [18:0] Wgt_1_48, // sfix19_En18 
  input [18:0] Wgt_1_49, // sfix19_En18 
  input [18:0] Wgt_1_50, // sfix19_En18 
  input [18:0] Wgt_1_51, // sfix19_En18 
  input [18:0] Wgt_1_52, // sfix19_En18 
  input [18:0] Wgt_1_53, // sfix19_En18 
  input [18:0] Wgt_1_54, // sfix19_En18 
  input [18:0] Wgt_1_55, // sfix19_En18 
  input [18:0] Wgt_1_56, // sfix19_En18 
  input [18:0] Wgt_1_57, // sfix19_En18 
  input [18:0] Wgt_1_58, // sfix19_En18 
  input [18:0] Wgt_1_59, // sfix19_En18 
  input [18:0] Wgt_1_60, // sfix19_En18 
  input [18:0] Wgt_1_61, // sfix19_En18 
  input [18:0] Wgt_1_62, // sfix19_En18 
  input [18:0] Wgt_1_63, // sfix19_En18 
  input [18:0] Wgt_1_64, // sfix19_En18 
  input [18:0] Wgt_1_65, // sfix19_En18 
  input [18:0] Wgt_1_66, // sfix19_En18 
  input [18:0] Wgt_1_67, // sfix19_En18 
  input [18:0] Wgt_1_68, // sfix19_En18 
  input [18:0] Wgt_1_69, // sfix19_En18 
  input [18:0] Wgt_1_70, // sfix19_En18 
  input [18:0] Wgt_1_71, // sfix19_En18 
  input [18:0] Wgt_1_72, // sfix19_En18 
  input [18:0] Wgt_1_73, // sfix19_En18 
  input [18:0] Wgt_1_74, // sfix19_En18 
  input [18:0] Wgt_1_75, // sfix19_En18 
  input [18:0] Wgt_1_76, // sfix19_En18 
  input [18:0] Wgt_1_77, // sfix19_En18 
  input [18:0] Wgt_1_78, // sfix19_En18 
  input [18:0] Wgt_1_79, // sfix19_En18 
  input [18:0] Wgt_1_80, // sfix19_En18 
  input [18:0] Wgt_1_81, // sfix19_En18 
  input [18:0] Wgt_1_82, // sfix19_En18 
  input [18:0] Wgt_1_83, // sfix19_En18 
  input [18:0] Wgt_1_84, // sfix19_En18 
  input [18:0] Wgt_1_85, // sfix19_En18 
  input [18:0] Wgt_1_86, // sfix19_En18 
  input [18:0] Wgt_1_87, // sfix19_En18 
  input [18:0] Wgt_1_88, // sfix19_En18 
  input [18:0] Wgt_1_89, // sfix19_En18 
  input [18:0] Wgt_1_90, // sfix19_En18 
  input [18:0] Wgt_1_91, // sfix19_En18 
  input [18:0] Wgt_1_92, // sfix19_En18 
  input [18:0] Wgt_1_93, // sfix19_En18 
  input [18:0] Wgt_1_94, // sfix19_En18 
  input [18:0] Wgt_1_95, // sfix19_En18 
  input [18:0] Wgt_1_96, // sfix19_En18 
  input [18:0] Wgt_1_97, // sfix19_En18 
  input [18:0] Wgt_1_98, // sfix19_En18 
  input [18:0] Wgt_1_99, // sfix19_En18 
  input [18:0] Wgt_1_100, // sfix19_En18 
  input [18:0] Wgt_1_101, // sfix19_En18 
  input [18:0] Wgt_1_102, // sfix19_En18 
  input [18:0] Wgt_1_103, // sfix19_En18 
  input [18:0] Wgt_1_104, // sfix19_En18 
  input [18:0] Wgt_1_105, // sfix19_En18 
  input [18:0] Wgt_1_106, // sfix19_En18 
  input [18:0] Wgt_1_107, // sfix19_En18 
  input [18:0] Wgt_1_108, // sfix19_En18 
  input [18:0] Wgt_1_109, // sfix19_En18 
  input [18:0] Wgt_1_110, // sfix19_En18 
  input [18:0] Wgt_1_111, // sfix19_En18 
  input [18:0] Wgt_1_112, // sfix19_En18 
  input [18:0] Wgt_1_113, // sfix19_En18 
  input [18:0] Wgt_1_114, // sfix19_En18 
  input [18:0] Wgt_1_115, // sfix19_En18 
  input [18:0] Wgt_1_116, // sfix19_En18 
  input [18:0] Wgt_1_117, // sfix19_En18 
  input [18:0] Wgt_1_118, // sfix19_En18 
  input [18:0] Wgt_1_119, // sfix19_En18 
  input [18:0] Wgt_1_120, // sfix19_En18 
  input [18:0] Wgt_1_121, // sfix19_En18 
  input [18:0] Wgt_1_122, // sfix19_En18 
  input [18:0] Wgt_1_123, // sfix19_En18 
  input [18:0] Wgt_1_124, // sfix19_En18 
  input [18:0] Wgt_1_125, // sfix19_En18 
  input [18:0] Wgt_1_126, // sfix19_En18 
  input [18:0] Wgt_1_127, // sfix19_En18 
  input [18:0] Wgt_1_128, // sfix19_En18 
  input [18:0] Wgt_1_129, // sfix19_En18 
  input [18:0] Wgt_1_130, // sfix19_En18 
  input [18:0] Wgt_1_131, // sfix19_En18 
  input [18:0] Wgt_1_132, // sfix19_En18 
  input [18:0] Wgt_1_133, // sfix19_En18 
  input [18:0] Wgt_1_134, // sfix19_En18 
  input [18:0] Wgt_1_135, // sfix19_En18 
  input [18:0] Wgt_1_136, // sfix19_En18 
  input [18:0] Wgt_1_137, // sfix19_En18 
  input [18:0] Wgt_1_138, // sfix19_En18 
  input [18:0] Wgt_1_139, // sfix19_En18 
  input [18:0] Wgt_1_140, // sfix19_En18 
  input [18:0] Wgt_1_141, // sfix19_En18 
  input [18:0] Wgt_1_142, // sfix19_En18 
  input [18:0] Wgt_1_143, // sfix19_En18 
  input [18:0] Wgt_1_144, // sfix19_En18 
  input [18:0] Wgt_1_145, // sfix19_En18 
  input [18:0] Wgt_1_146, // sfix19_En18 
  input [18:0] Wgt_1_147, // sfix19_En18 
  input [18:0] Wgt_1_148, // sfix19_En18 
  input [18:0] Wgt_1_149, // sfix19_En18 
  input [18:0] Wgt_1_150, // sfix19_En18 
  input [18:0] Wgt_1_151, // sfix19_En18 
  input [18:0] Wgt_1_152, // sfix19_En18 
  input [18:0] Wgt_1_153, // sfix19_En18 
  input [18:0] Wgt_1_154, // sfix19_En18 
  input [18:0] Wgt_1_155, // sfix19_En18 
  input [18:0] Wgt_1_156, // sfix19_En18 
  input [18:0] Wgt_1_157, // sfix19_En18 
  input [18:0] Wgt_1_158, // sfix19_En18 
  input [18:0] Wgt_1_159, // sfix19_En18 
  input [18:0] Wgt_1_160, // sfix19_En18 
  input [18:0] Wgt_1_161, // sfix19_En18 
  input [18:0] Wgt_1_162, // sfix19_En18 
  input [18:0] Wgt_1_163, // sfix19_En18 
  input [18:0] Wgt_1_164, // sfix19_En18 
  input [18:0] Wgt_1_165, // sfix19_En18 
  input [18:0] Wgt_1_166, // sfix19_En18 
  input [18:0] Wgt_1_167, // sfix19_En18 
  input [18:0] Wgt_1_168, // sfix19_En18 
  input [18:0] Wgt_1_169, // sfix19_En18 
  input [18:0] Wgt_1_170, // sfix19_En18 
  input [18:0] Wgt_1_171, // sfix19_En18 
  input [18:0] Wgt_1_172, // sfix19_En18 
  input [18:0] Wgt_1_173, // sfix19_En18 
  input [18:0] Wgt_1_174, // sfix19_En18 
  input [18:0] Wgt_1_175, // sfix19_En18 
  input [18:0] Wgt_1_176, // sfix19_En18 
  input [18:0] Wgt_1_177, // sfix19_En18 
  input [18:0] Wgt_1_178, // sfix19_En18 
  input [18:0] Wgt_1_179, // sfix19_En18 
  input [18:0] Wgt_1_180, // sfix19_En18 
  input [18:0] Wgt_1_181, // sfix19_En18 
  input [18:0] Wgt_1_182, // sfix19_En18 
  input [18:0] Wgt_1_183, // sfix19_En18 
  input [18:0] Wgt_1_184, // sfix19_En18 
  input [18:0] Wgt_1_185, // sfix19_En18 
  input [18:0] Wgt_1_186, // sfix19_En18 
  input [18:0] Wgt_1_187, // sfix19_En18 
  input [18:0] Wgt_1_188, // sfix19_En18 
  input [18:0] Wgt_1_189, // sfix19_En18 
  input [18:0] Wgt_1_190, // sfix19_En18 
  input [18:0] Wgt_1_191, // sfix19_En18 
  input [18:0] Wgt_1_192, // sfix19_En18 
  input [18:0] Wgt_1_193, // sfix19_En18 
  input [18:0] Wgt_1_194, // sfix19_En18 
  input [18:0] Wgt_1_195, // sfix19_En18 
  input [18:0] Wgt_1_196, // sfix19_En18 
  input [18:0] Wgt_1_197, // sfix19_En18 
  input [18:0] Wgt_1_198, // sfix19_En18 
  input [18:0] Wgt_1_199, // sfix19_En18 
  input [18:0] Wgt_1_200, // sfix19_En18 
  input [18:0] Wgt_1_201, // sfix19_En18 
  input [18:0] Wgt_1_202, // sfix19_En18 
  input [18:0] Wgt_1_203, // sfix19_En18 
  input [18:0] Wgt_1_204, // sfix19_En18 
  input [18:0] Wgt_1_205, // sfix19_En18 
  input [18:0] Wgt_1_206, // sfix19_En18 
  input [18:0] Wgt_1_207, // sfix19_En18 
  input [18:0] Wgt_1_208, // sfix19_En18 
  input [18:0] Wgt_1_209, // sfix19_En18 
  input [18:0] Wgt_1_210, // sfix19_En18 
  input [18:0] Wgt_1_211, // sfix19_En18 
  input [18:0] Wgt_1_212, // sfix19_En18 
  input [18:0] Wgt_1_213, // sfix19_En18 
  input [18:0] Wgt_1_214, // sfix19_En18 
  input [18:0] Wgt_1_215, // sfix19_En18 
  input [18:0] Wgt_1_216, // sfix19_En18 
  input [18:0] Wgt_1_217, // sfix19_En18 
  input [18:0] Wgt_1_218, // sfix19_En18 
  input [18:0] Wgt_1_219, // sfix19_En18 
  input [18:0] Wgt_1_220, // sfix19_En18 
  input [18:0] Wgt_1_221, // sfix19_En18 
  input [18:0] Wgt_1_222, // sfix19_En18 
  input [18:0] Wgt_1_223, // sfix19_En18 
  input [18:0] Wgt_1_224, // sfix19_En18 
  input [18:0] Wgt_1_225, // sfix19_En18 
  input [18:0] Wgt_1_226, // sfix19_En18 
  input [18:0] Wgt_1_227, // sfix19_En18 
  input [18:0] Wgt_1_228, // sfix19_En18 
  input [18:0] Wgt_1_229, // sfix19_En18 
  input [18:0] Wgt_1_230, // sfix19_En18 
  input [18:0] Wgt_1_231, // sfix19_En18 
  input [18:0] Wgt_1_232, // sfix19_En18 
  input [18:0] Wgt_1_233, // sfix19_En18 
  input [18:0] Wgt_1_234, // sfix19_En18 
  input [18:0] Wgt_1_235, // sfix19_En18 
  input [18:0] Wgt_1_236, // sfix19_En18 
  input [18:0] Wgt_1_237, // sfix19_En18 
  input [18:0] Wgt_1_238, // sfix19_En18 
  input [18:0] Wgt_1_239, // sfix19_En18 
  input [18:0] Wgt_1_240, // sfix19_En18 
  input [18:0] Wgt_1_241, // sfix19_En18 
  input [18:0] Wgt_1_242, // sfix19_En18 
  input [18:0] Wgt_1_243, // sfix19_En18 
  input [18:0] Wgt_1_244, // sfix19_En18 
  input [18:0] Wgt_1_245, // sfix19_En18 
  input [18:0] Wgt_1_246, // sfix19_En18 
  input [18:0] Wgt_1_247, // sfix19_En18 
  input [18:0] Wgt_1_248, // sfix19_En18 
  input [18:0] Wgt_1_249, // sfix19_En18 
  input [18:0] Wgt_1_250, // sfix19_En18 
  input [18:0] Wgt_1_251, // sfix19_En18 
  input [18:0] Wgt_1_252, // sfix19_En18 
  input [18:0] Wgt_1_253, // sfix19_En18 
  input [18:0] Wgt_1_254, // sfix19_En18 
  input [18:0] Wgt_1_255, // sfix19_En18 
  input [18:0] Wgt_1_256, // sfix19_En18 
  input [18:0] Wgt_1_257, // sfix19_En18 
  input [18:0] Wgt_1_258, // sfix19_En18 
  input [18:0] Wgt_1_259, // sfix19_En18 
  input [18:0] Wgt_1_260, // sfix19_En18 
  input [18:0] Wgt_1_261, // sfix19_En18 
  input [18:0] Wgt_1_262, // sfix19_En18 
  input [18:0] Wgt_1_263, // sfix19_En18 
  input [18:0] Wgt_1_264, // sfix19_En18 
  input [18:0] Wgt_1_265, // sfix19_En18 
  input [18:0] Wgt_1_266, // sfix19_En18 
  input [18:0] Wgt_1_267, // sfix19_En18 
  input [18:0] Wgt_1_268, // sfix19_En18 
  input [18:0] Wgt_1_269, // sfix19_En18 
  input [18:0] Wgt_1_270, // sfix19_En18 
  input [18:0] Wgt_1_271, // sfix19_En18 
  input [18:0] Wgt_1_272, // sfix19_En18 
  input [18:0] Wgt_1_273, // sfix19_En18 
  input [18:0] Wgt_1_274, // sfix19_En18 
  input [18:0] Wgt_1_275, // sfix19_En18 
  input [18:0] Wgt_1_276, // sfix19_En18 
  input [18:0] Wgt_1_277, // sfix19_En18 
  input [18:0] Wgt_1_278, // sfix19_En18 
  input [18:0] Wgt_1_279, // sfix19_En18 
  input [18:0] Wgt_1_280, // sfix19_En18 
  input [18:0] Wgt_1_281, // sfix19_En18 
  input [18:0] Wgt_1_282, // sfix19_En18 
  input [18:0] Wgt_1_283, // sfix19_En18 
  input [18:0] Wgt_1_284, // sfix19_En18 
  input [18:0] Wgt_1_285, // sfix19_En18 
  input [18:0] Wgt_1_286, // sfix19_En18 
  input [18:0] Wgt_1_287, // sfix19_En18 
  input [18:0] Wgt_1_288, // sfix19_En18 
  input [18:0] Wgt_1_289, // sfix19_En18 
  input [18:0] Wgt_1_290, // sfix19_En18 
  input [18:0] Wgt_1_291, // sfix19_En18 
  input [18:0] Wgt_1_292, // sfix19_En18 
  input [18:0] Wgt_1_293, // sfix19_En18 
  input [18:0] Wgt_1_294, // sfix19_En18 
  input [18:0] Wgt_1_295, // sfix19_En18 
  input [18:0] Wgt_1_296, // sfix19_En18 
  input [18:0] Wgt_1_297, // sfix19_En18 
  input [18:0] Wgt_1_298, // sfix19_En18 
  input [18:0] Wgt_1_299, // sfix19_En18 
  input [18:0] Wgt_1_300, // sfix19_En18 
  input [18:0] Wgt_1_301, // sfix19_En18 
  input [18:0] Wgt_1_302, // sfix19_En18 
  input [18:0] Wgt_1_303, // sfix19_En18 
  input [18:0] Wgt_1_304, // sfix19_En18 
  input [18:0] Wgt_1_305, // sfix19_En18 
  input [18:0] Wgt_1_306, // sfix19_En18 
  input [18:0] Wgt_1_307, // sfix19_En18 
  input [18:0] Wgt_1_308, // sfix19_En18 
  input [18:0] Wgt_1_309, // sfix19_En18 
  input [18:0] Wgt_1_310, // sfix19_En18 
  input [18:0] Wgt_1_311, // sfix19_En18 
  input [18:0] Wgt_1_312, // sfix19_En18 
  input [18:0] Wgt_1_313, // sfix19_En18 
  input [18:0] Wgt_1_314, // sfix19_En18 
  input [18:0] Wgt_1_315, // sfix19_En18 
  input [18:0] Wgt_1_316, // sfix19_En18 
  input [18:0] Wgt_1_317, // sfix19_En18 
  input [18:0] Wgt_1_318, // sfix19_En18 
  input [18:0] Wgt_1_319, // sfix19_En18 
  input [18:0] Wgt_1_320, // sfix19_En18 
  input [18:0] Wgt_1_321, // sfix19_En18 
  input [18:0] Wgt_1_322, // sfix19_En18 
  input [18:0] Wgt_1_323, // sfix19_En18 
  input [18:0] Wgt_1_324, // sfix19_En18 
  input [18:0] Wgt_1_325, // sfix19_En18 
  input [18:0] Wgt_1_326, // sfix19_En18 
  input [18:0] Wgt_1_327, // sfix19_En18 
  input [18:0] Wgt_1_328, // sfix19_En18 
  input [18:0] Wgt_1_329, // sfix19_En18 
  input [18:0] Wgt_1_330, // sfix19_En18 
  input [18:0] Wgt_1_331, // sfix19_En18 
  input [18:0] Wgt_1_332, // sfix19_En18 
  input [18:0] Wgt_1_333, // sfix19_En18 
  input [18:0] Wgt_1_334, // sfix19_En18 
  input [18:0] Wgt_1_335, // sfix19_En18 
  input [18:0] Wgt_1_336, // sfix19_En18 
  input [18:0] Wgt_1_337, // sfix19_En18 
  input [18:0] Wgt_1_338, // sfix19_En18 
  input [18:0] Wgt_1_339, // sfix19_En18 
  input [18:0] Wgt_1_340, // sfix19_En18 
  input [18:0] Wgt_1_341, // sfix19_En18 
  input [18:0] Wgt_1_342, // sfix19_En18 
  input [18:0] Wgt_1_343, // sfix19_En18 
  input [18:0] Wgt_1_344, // sfix19_En18 
  input [18:0] Wgt_1_345, // sfix19_En18 
  input [18:0] Wgt_1_346, // sfix19_En18 
  input [18:0] Wgt_1_347, // sfix19_En18 
  input [18:0] Wgt_1_348, // sfix19_En18 
  input [18:0] Wgt_1_349, // sfix19_En18 
  input [18:0] Wgt_1_350, // sfix19_En18 
  input [18:0] Wgt_1_351, // sfix19_En18 
  input [18:0] Wgt_1_352, // sfix19_En18 
  input [18:0] Wgt_1_353, // sfix19_En18 
  input [18:0] Wgt_1_354, // sfix19_En18 
  input [18:0] Wgt_1_355, // sfix19_En18 
  input [18:0] Wgt_1_356, // sfix19_En18 
  input [18:0] Wgt_1_357, // sfix19_En18 
  input [18:0] Wgt_1_358, // sfix19_En18 
  input [18:0] Wgt_1_359, // sfix19_En18 
  input [18:0] Wgt_1_360, // sfix19_En18 
  input [18:0] Wgt_1_361, // sfix19_En18 
  input [18:0] Wgt_1_362, // sfix19_En18 
  input [18:0] Wgt_1_363, // sfix19_En18 
  input [18:0] Wgt_1_364, // sfix19_En18 
  input [18:0] Wgt_1_365, // sfix19_En18 
  input [18:0] Wgt_1_366, // sfix19_En18 
  input [18:0] Wgt_1_367, // sfix19_En18 
  input [18:0] Wgt_1_368, // sfix19_En18 
  input [18:0] Wgt_1_369, // sfix19_En18 
  input [18:0] Wgt_1_370, // sfix19_En18 
  input [18:0] Wgt_1_371, // sfix19_En18 
  input [18:0] Wgt_1_372, // sfix19_En18 
  input [18:0] Wgt_1_373, // sfix19_En18 
  input [18:0] Wgt_1_374, // sfix19_En18 
  input [18:0] Wgt_1_375, // sfix19_En18 
  input [18:0] Wgt_1_376, // sfix19_En18 
  input [18:0] Wgt_1_377, // sfix19_En18 
  input [18:0] Wgt_1_378, // sfix19_En18 
  input [18:0] Wgt_1_379, // sfix19_En18 
  input [18:0] Wgt_1_380, // sfix19_En18 
  input [18:0] Wgt_1_381, // sfix19_En18 
  input [18:0] Wgt_1_382, // sfix19_En18 
  input [18:0] Wgt_1_383, // sfix19_En18 
  input [18:0] Wgt_1_384, // sfix19_En18 
  input [18:0] Wgt_1_385, // sfix19_En18 
  input [18:0] Wgt_1_386, // sfix19_En18 
  input [18:0] Wgt_1_387, // sfix19_En18 
  input [18:0] Wgt_1_388, // sfix19_En18 
  input [18:0] Wgt_1_389, // sfix19_En18 
  input [18:0] Wgt_1_390, // sfix19_En18 
  input [18:0] Wgt_1_391, // sfix19_En18 
  input [18:0] Wgt_1_392, // sfix19_En18 
  input [18:0] Wgt_1_393, // sfix19_En18 
  input [18:0] Wgt_1_394, // sfix19_En18 
  input [18:0] Wgt_1_395, // sfix19_En18 
  input [18:0] Wgt_1_396, // sfix19_En18 
  input [18:0] Wgt_1_397, // sfix19_En18 
  input [18:0] Wgt_1_398, // sfix19_En18 
  input [18:0] Wgt_1_399, // sfix19_En18 
  input [18:0] Wgt_1_400, // sfix19_En18 
  input [18:0] Wgt_1_401, // sfix19_En18 
  input [18:0] Wgt_1_402, // sfix19_En18 
  input [18:0] Wgt_1_403, // sfix19_En18 
  input [18:0] Wgt_1_404, // sfix19_En18 
  input [18:0] Wgt_1_405, // sfix19_En18 
  input [18:0] Wgt_1_406, // sfix19_En18 
  input [18:0] Wgt_1_407, // sfix19_En18 
  input [18:0] Wgt_1_408, // sfix19_En18 
  input [18:0] Wgt_1_409, // sfix19_En18 
  input [18:0] Wgt_1_410, // sfix19_En18 
  input [18:0] Wgt_1_411, // sfix19_En18 
  input [18:0] Wgt_1_412, // sfix19_En18 
  input [18:0] Wgt_1_413, // sfix19_En18 
  input [18:0] Wgt_1_414, // sfix19_En18 
  input [18:0] Wgt_1_415, // sfix19_En18 
  input [18:0] Wgt_1_416, // sfix19_En18 
  input [18:0] Wgt_1_417, // sfix19_En18 
  input [18:0] Wgt_1_418, // sfix19_En18 
  input [18:0] Wgt_1_419, // sfix19_En18 
  input [18:0] Wgt_1_420, // sfix19_En18 
  input [18:0] Wgt_1_421, // sfix19_En18 
  input [18:0] Wgt_1_422, // sfix19_En18 
  input [18:0] Wgt_1_423, // sfix19_En18 
  input [18:0] Wgt_1_424, // sfix19_En18 
  input [18:0] Wgt_1_425, // sfix19_En18 
  input [18:0] Wgt_1_426, // sfix19_En18 
  input [18:0] Wgt_1_427, // sfix19_En18 
  input [18:0] Wgt_1_428, // sfix19_En18 
  input [18:0] Wgt_1_429, // sfix19_En18 
  input [18:0] Wgt_1_430, // sfix19_En18 
  input [18:0] Wgt_1_431, // sfix19_En18 
  input [18:0] Wgt_1_432, // sfix19_En18 
  input [18:0] Wgt_1_433, // sfix19_En18 
  input [18:0] Wgt_1_434, // sfix19_En18 
  input [18:0] Wgt_1_435, // sfix19_En18 
  input [18:0] Wgt_1_436, // sfix19_En18 
  input [18:0] Wgt_1_437, // sfix19_En18 
  input [18:0] Wgt_1_438, // sfix19_En18 
  input [18:0] Wgt_1_439, // sfix19_En18 
  input [18:0] Wgt_1_440, // sfix19_En18 
  input [18:0] Wgt_1_441, // sfix19_En18 
  input [18:0] Wgt_1_442, // sfix19_En18 
  input [18:0] Wgt_1_443, // sfix19_En18 
  input [18:0] Wgt_1_444, // sfix19_En18 
  input [18:0] Wgt_1_445, // sfix19_En18 
  input [18:0] Wgt_1_446, // sfix19_En18 
  input [18:0] Wgt_1_447, // sfix19_En18 
  input [18:0] Wgt_1_448, // sfix19_En18 
  input [18:0] Wgt_1_449, // sfix19_En18 
  input [18:0] Wgt_1_450, // sfix19_En18 
  input [18:0] Wgt_1_451, // sfix19_En18 
  input [18:0] Wgt_1_452, // sfix19_En18 
  input [18:0] Wgt_1_453, // sfix19_En18 
  input [18:0] Wgt_1_454, // sfix19_En18 
  input [18:0] Wgt_1_455, // sfix19_En18 
  input [18:0] Wgt_1_456, // sfix19_En18 
  input [18:0] Wgt_1_457, // sfix19_En18 
  input [18:0] Wgt_1_458, // sfix19_En18 
  input [18:0] Wgt_1_459, // sfix19_En18 
  input [18:0] Wgt_1_460, // sfix19_En18 
  input [18:0] Wgt_1_461, // sfix19_En18 
  input [18:0] Wgt_1_462, // sfix19_En18 
  input [18:0] Wgt_1_463, // sfix19_En18 
  input [18:0] Wgt_1_464, // sfix19_En18 
  input [18:0] Wgt_1_465, // sfix19_En18 
  input [18:0] Wgt_1_466, // sfix19_En18 
  input [18:0] Wgt_1_467, // sfix19_En18 
  input [18:0] Wgt_1_468, // sfix19_En18 
  input [18:0] Wgt_1_469, // sfix19_En18 
  input [18:0] Wgt_1_470, // sfix19_En18 
  input [18:0] Wgt_1_471, // sfix19_En18 
  input [18:0] Wgt_1_472, // sfix19_En18 
  input [18:0] Wgt_1_473, // sfix19_En18 
  input [18:0] Wgt_1_474, // sfix19_En18 
  input [18:0] Wgt_1_475, // sfix19_En18 
  input [18:0] Wgt_1_476, // sfix19_En18 
  input [18:0] Wgt_1_477, // sfix19_En18 
  input [18:0] Wgt_1_478, // sfix19_En18 
  input [18:0] Wgt_1_479, // sfix19_En18 
  input [18:0] Wgt_1_480, // sfix19_En18 
  input [18:0] Wgt_1_481, // sfix19_En18 
  input [18:0] Wgt_1_482, // sfix19_En18 
  input [18:0] Wgt_1_483, // sfix19_En18 
  input [18:0] Wgt_1_484, // sfix19_En18 
  input [18:0] Wgt_1_485, // sfix19_En18 
  input [18:0] Wgt_1_486, // sfix19_En18 
  input [18:0] Wgt_1_487, // sfix19_En18 
  input [18:0] Wgt_1_488, // sfix19_En18 
  input [18:0] Wgt_1_489, // sfix19_En18 
  input [18:0] Wgt_1_490, // sfix19_En18 
  input [18:0] Wgt_1_491, // sfix19_En18 
  input [18:0] Wgt_1_492, // sfix19_En18 
  input [18:0] Wgt_1_493, // sfix19_En18 
  input [18:0] Wgt_1_494, // sfix19_En18 
  input [18:0] Wgt_1_495, // sfix19_En18 
  input [18:0] Wgt_1_496, // sfix19_En18 
  input [18:0] Wgt_1_497, // sfix19_En18 
  input [18:0] Wgt_1_498, // sfix19_En18 
  input [18:0] Wgt_1_499, // sfix19_En18 
  input [18:0] Wgt_1_500, // sfix19_En18 
  input [18:0] Wgt_1_501, // sfix19_En18 
  input [18:0] Wgt_1_502, // sfix19_En18 
  input [18:0] Wgt_1_503, // sfix19_En18 
  input [18:0] Wgt_1_504, // sfix19_En18 
  input [18:0] Wgt_1_505, // sfix19_En18 
  input [18:0] Wgt_1_506, // sfix19_En18 
  input [18:0] Wgt_1_507, // sfix19_En18 
  input [18:0] Wgt_1_508, // sfix19_En18 
  input [18:0] Wgt_1_509, // sfix19_En18 
  input [18:0] Wgt_1_510, // sfix19_En18 
  input [18:0] Wgt_1_511, // sfix19_En18 
  input [18:0] Wgt_1_512, // sfix19_En18 
  input [18:0] Wgt_1_513, // sfix19_En18 
  input [18:0] Wgt_1_514, // sfix19_En18 
  input [18:0] Wgt_1_515, // sfix19_En18 
  input [18:0] Wgt_1_516, // sfix19_En18 
  input [18:0] Wgt_1_517, // sfix19_En18 
  input [18:0] Wgt_1_518, // sfix19_En18 
  input [18:0] Wgt_1_519, // sfix19_En18 
  input [18:0] Wgt_1_520, // sfix19_En18 
  input [18:0] Wgt_1_521, // sfix19_En18 
  input [18:0] Wgt_1_522, // sfix19_En18 
  input [18:0] Wgt_1_523, // sfix19_En18 
  input [18:0] Wgt_1_524, // sfix19_En18 
  input [18:0] Wgt_1_525, // sfix19_En18 
  input [18:0] Wgt_1_526, // sfix19_En18 
  input [18:0] Wgt_1_527, // sfix19_En18 
  input [18:0] Wgt_1_528, // sfix19_En18 
  input [18:0] Wgt_1_529, // sfix19_En18 
  input [18:0] Wgt_1_530, // sfix19_En18 
  input [18:0] Wgt_1_531, // sfix19_En18 
  input [18:0] Wgt_1_532, // sfix19_En18 
  input [18:0] Wgt_1_533, // sfix19_En18 
  input [18:0] Wgt_1_534, // sfix19_En18 
  input [18:0] Wgt_1_535, // sfix19_En18 
  input [18:0] Wgt_1_536, // sfix19_En18 
  input [18:0] Wgt_1_537, // sfix19_En18 
  input [18:0] Wgt_1_538, // sfix19_En18 
  input [18:0] Wgt_1_539, // sfix19_En18 
  input [18:0] Wgt_1_540, // sfix19_En18 
  input [18:0] Wgt_1_541, // sfix19_En18 
  input [18:0] Wgt_1_542, // sfix19_En18 
  input [18:0] Wgt_1_543, // sfix19_En18 
  input [18:0] Wgt_1_544, // sfix19_En18 
  input [18:0] Wgt_1_545, // sfix19_En18 
  input [18:0] Wgt_1_546, // sfix19_En18 
  input [18:0] Wgt_1_547, // sfix19_En18 
  input [18:0] Wgt_1_548, // sfix19_En18 
  input [18:0] Wgt_1_549, // sfix19_En18 
  input [18:0] Wgt_1_550, // sfix19_En18 
  input [18:0] Wgt_1_551, // sfix19_En18 
  input [18:0] Wgt_1_552, // sfix19_En18 
  input [18:0] Wgt_1_553, // sfix19_En18 
  input [18:0] Wgt_1_554, // sfix19_En18 
  input [18:0] Wgt_1_555, // sfix19_En18 
  input [18:0] Wgt_1_556, // sfix19_En18 
  input [18:0] Wgt_1_557, // sfix19_En18 
  input [18:0] Wgt_1_558, // sfix19_En18 
  input [18:0] Wgt_1_559, // sfix19_En18 
  input [18:0] Wgt_1_560, // sfix19_En18 
  input [18:0] Wgt_1_561, // sfix19_En18 
  input [18:0] Wgt_1_562, // sfix19_En18 
  input [18:0] Wgt_1_563, // sfix19_En18 
  input [18:0] Wgt_1_564, // sfix19_En18 
  input [18:0] Wgt_1_565, // sfix19_En18 
  input [18:0] Wgt_1_566, // sfix19_En18 
  input [18:0] Wgt_1_567, // sfix19_En18 
  input [18:0] Wgt_1_568, // sfix19_En18 
  input [18:0] Wgt_1_569, // sfix19_En18 
  input [18:0] Wgt_1_570, // sfix19_En18 
  input [18:0] Wgt_1_571, // sfix19_En18 
  input [18:0] Wgt_1_572, // sfix19_En18 
  input [18:0] Wgt_1_573, // sfix19_En18 
  input [18:0] Wgt_1_574, // sfix19_En18 
  input [18:0] Wgt_1_575, // sfix19_En18 
  input [18:0] Wgt_1_576, // sfix19_En18 
  input [18:0] Wgt_1_577, // sfix19_En18 
  input [18:0] Wgt_1_578, // sfix19_En18 
  input [18:0] Wgt_1_579, // sfix19_En18 
  input [18:0] Wgt_1_580, // sfix19_En18 
  input [18:0] Wgt_1_581, // sfix19_En18 
  input [18:0] Wgt_1_582, // sfix19_En18 
  input [18:0] Wgt_1_583, // sfix19_En18 
  input [18:0] Wgt_1_584, // sfix19_En18 
  input [18:0] Wgt_1_585, // sfix19_En18 
  input [18:0] Wgt_1_586, // sfix19_En18 
  input [18:0] Wgt_1_587, // sfix19_En18 
  input [18:0] Wgt_1_588, // sfix19_En18 
  input [18:0] Wgt_1_589, // sfix19_En18 
  input [18:0] Wgt_1_590, // sfix19_En18 
  input [18:0] Wgt_1_591, // sfix19_En18 
  input [18:0] Wgt_1_592, // sfix19_En18 
  input [18:0] Wgt_1_593, // sfix19_En18 
  input [18:0] Wgt_1_594, // sfix19_En18 
  input [18:0] Wgt_1_595, // sfix19_En18 
  input [18:0] Wgt_1_596, // sfix19_En18 
  input [18:0] Wgt_1_597, // sfix19_En18 
  input [18:0] Wgt_1_598, // sfix19_En18 
  input [18:0] Wgt_1_599, // sfix19_En18 
  input [18:0] Wgt_1_600, // sfix19_En18 
  input [18:0] Wgt_1_601, // sfix19_En18 
  input [18:0] Wgt_1_602, // sfix19_En18 
  input [18:0] Wgt_1_603, // sfix19_En18 
  input [18:0] Wgt_1_604, // sfix19_En18 
  input [18:0] Wgt_1_605, // sfix19_En18 
  input [18:0] Wgt_1_606, // sfix19_En18 
  input [18:0] Wgt_1_607, // sfix19_En18 
  input [18:0] Wgt_1_608, // sfix19_En18 
  input [18:0] Wgt_1_609, // sfix19_En18 
  input [18:0] Wgt_1_610, // sfix19_En18 
  input [18:0] Wgt_1_611, // sfix19_En18 
  input [18:0] Wgt_1_612, // sfix19_En18 
  input [18:0] Wgt_1_613, // sfix19_En18 
  input [18:0] Wgt_1_614, // sfix19_En18 
  input [18:0] Wgt_1_615, // sfix19_En18 
  input [18:0] Wgt_1_616, // sfix19_En18 
  input [18:0] Wgt_1_617, // sfix19_En18 
  input [18:0] Wgt_1_618, // sfix19_En18 
  input [18:0] Wgt_1_619, // sfix19_En18 
  input [18:0] Wgt_1_620, // sfix19_En18 
  input [18:0] Wgt_1_621, // sfix19_En18 
  input [18:0] Wgt_1_622, // sfix19_En18 
  input [18:0] Wgt_1_623, // sfix19_En18 
  input [18:0] Wgt_1_624, // sfix19_En18 
  input [18:0] Wgt_1_625, // sfix19_En18 
  input [18:0] Wgt_1_626, // sfix19_En18 
  input [18:0] Wgt_1_627, // sfix19_En18 
  input [18:0] Wgt_1_628, // sfix19_En18 
  input [18:0] Wgt_1_629, // sfix19_En18 
  input [18:0] Wgt_1_630, // sfix19_En18 
  input [18:0] Wgt_1_631, // sfix19_En18 
  input [18:0] Wgt_1_632, // sfix19_En18 
  input [18:0] Wgt_1_633, // sfix19_En18 
  input [18:0] Wgt_1_634, // sfix19_En18 
  input [18:0] Wgt_1_635, // sfix19_En18 
  input [18:0] Wgt_1_636, // sfix19_En18 
  input [18:0] Wgt_1_637, // sfix19_En18 
  input [18:0] Wgt_1_638, // sfix19_En18 
  input [18:0] Wgt_1_639, // sfix19_En18 
  input [18:0] Wgt_1_640, // sfix19_En18 
  input [18:0] Wgt_1_641, // sfix19_En18 
  input [18:0] Wgt_1_642, // sfix19_En18 
  input [18:0] Wgt_1_643, // sfix19_En18 
  input [18:0] Wgt_1_644, // sfix19_En18 
  input [18:0] Wgt_1_645, // sfix19_En18 
  input [18:0] Wgt_1_646, // sfix19_En18 
  input [18:0] Wgt_1_647, // sfix19_En18 
  input [18:0] Wgt_1_648, // sfix19_En18 
  input [18:0] Wgt_1_649, // sfix19_En18 
  input [18:0] Wgt_1_650, // sfix19_En18 
  input [18:0] Wgt_1_651, // sfix19_En18 
  input [18:0] Wgt_1_652, // sfix19_En18 
  input [18:0] Wgt_1_653, // sfix19_En18 
  input [18:0] Wgt_1_654, // sfix19_En18 
  input [18:0] Wgt_1_655, // sfix19_En18 
  input [18:0] Wgt_1_656, // sfix19_En18 
  input [18:0] Wgt_1_657, // sfix19_En18 
  input [18:0] Wgt_1_658, // sfix19_En18 
  input [18:0] Wgt_1_659, // sfix19_En18 
  input [18:0] Wgt_1_660, // sfix19_En18 
  input [18:0] Wgt_1_661, // sfix19_En18 
  input [18:0] Wgt_1_662, // sfix19_En18 
  input [18:0] Wgt_1_663, // sfix19_En18 
  input [18:0] Wgt_1_664, // sfix19_En18 
  input [18:0] Wgt_1_665, // sfix19_En18 
  input [18:0] Wgt_1_666, // sfix19_En18 
  input [18:0] Wgt_1_667, // sfix19_En18 
  input [18:0] Wgt_1_668, // sfix19_En18 
  input [18:0] Wgt_1_669, // sfix19_En18 
  input [18:0] Wgt_1_670, // sfix19_En18 
  input [18:0] Wgt_1_671, // sfix19_En18 
  input [18:0] Wgt_1_672, // sfix19_En18 
  input [18:0] Wgt_1_673, // sfix19_En18 
  input [18:0] Wgt_1_674, // sfix19_En18 
  input [18:0] Wgt_1_675, // sfix19_En18 
  input [18:0] Wgt_1_676, // sfix19_En18 
  input [18:0] Wgt_1_677, // sfix19_En18 
  input [18:0] Wgt_1_678, // sfix19_En18 
  input [18:0] Wgt_1_679, // sfix19_En18 
  input [18:0] Wgt_1_680, // sfix19_En18 
  input [18:0] Wgt_1_681, // sfix19_En18 
  input [18:0] Wgt_1_682, // sfix19_En18 
  input [18:0] Wgt_1_683, // sfix19_En18 
  input [18:0] Wgt_1_684, // sfix19_En18 
  input [18:0] Wgt_1_685, // sfix19_En18 
  input [18:0] Wgt_1_686, // sfix19_En18 
  input [18:0] Wgt_1_687, // sfix19_En18 
  input [18:0] Wgt_1_688, // sfix19_En18 
  input [18:0] Wgt_1_689, // sfix19_En18 
  input [18:0] Wgt_1_690, // sfix19_En18 
  input [18:0] Wgt_1_691, // sfix19_En18 
  input [18:0] Wgt_1_692, // sfix19_En18 
  input [18:0] Wgt_1_693, // sfix19_En18 
  input [18:0] Wgt_1_694, // sfix19_En18 
  input [18:0] Wgt_1_695, // sfix19_En18 
  input [18:0] Wgt_1_696, // sfix19_En18 
  input [18:0] Wgt_1_697, // sfix19_En18 
  input [18:0] Wgt_1_698, // sfix19_En18 
  input [18:0] Wgt_1_699, // sfix19_En18 
  input [18:0] Wgt_1_700, // sfix19_En18 
  input [18:0] Wgt_1_701, // sfix19_En18 
  input [18:0] Wgt_1_702, // sfix19_En18 
  input [18:0] Wgt_1_703, // sfix19_En18 
  input [18:0] Wgt_1_704, // sfix19_En18 
  input [18:0] Wgt_1_705, // sfix19_En18 
  input [18:0] Wgt_1_706, // sfix19_En18 
  input [18:0] Wgt_1_707, // sfix19_En18 
  input [18:0] Wgt_1_708, // sfix19_En18 
  input [18:0] Wgt_1_709, // sfix19_En18 
  input [18:0] Wgt_1_710, // sfix19_En18 
  input [18:0] Wgt_1_711, // sfix19_En18 
  input [18:0] Wgt_1_712, // sfix19_En18 
  input [18:0] Wgt_1_713, // sfix19_En18 
  input [18:0] Wgt_1_714, // sfix19_En18 
  input [18:0] Wgt_1_715, // sfix19_En18 
  input [18:0] Wgt_1_716, // sfix19_En18 
  input [18:0] Wgt_1_717, // sfix19_En18 
  input [18:0] Wgt_1_718, // sfix19_En18 
  input [18:0] Wgt_1_719, // sfix19_En18 
  input [18:0] Wgt_1_720, // sfix19_En18 
  input [18:0] Wgt_1_721, // sfix19_En18 
  input [18:0] Wgt_1_722, // sfix19_En18 
  input [18:0] Wgt_1_723, // sfix19_En18 
  input [18:0] Wgt_1_724, // sfix19_En18 
  input [18:0] Wgt_1_725, // sfix19_En18 
  input [18:0] Wgt_1_726, // sfix19_En18 
  input [18:0] Wgt_1_727, // sfix19_En18 
  input [18:0] Wgt_1_728, // sfix19_En18 
  input [18:0] Wgt_1_729, // sfix19_En18 
  input [18:0] Wgt_1_730, // sfix19_En18 
  input [18:0] Wgt_1_731, // sfix19_En18 
  input [18:0] Wgt_1_732, // sfix19_En18 
  input [18:0] Wgt_1_733, // sfix19_En18 
  input [18:0] Wgt_1_734, // sfix19_En18 
  input [18:0] Wgt_1_735, // sfix19_En18 
  input [18:0] Wgt_1_736, // sfix19_En18 
  input [18:0] Wgt_1_737, // sfix19_En18 
  input [18:0] Wgt_1_738, // sfix19_En18 
  input [18:0] Wgt_1_739, // sfix19_En18 
  input [18:0] Wgt_1_740, // sfix19_En18 
  input [18:0] Wgt_1_741, // sfix19_En18 
  input [18:0] Wgt_1_742, // sfix19_En18 
  input [18:0] Wgt_1_743, // sfix19_En18 
  input [18:0] Wgt_1_744, // sfix19_En18 
  input [18:0] Wgt_1_745, // sfix19_En18 
  input [18:0] Wgt_1_746, // sfix19_En18 
  input [18:0] Wgt_1_747, // sfix19_En18 
  input [18:0] Wgt_1_748, // sfix19_En18 
  input [18:0] Wgt_1_749, // sfix19_En18 
  input [18:0] Wgt_1_750, // sfix19_En18 
  input [18:0] Wgt_1_751, // sfix19_En18 
  input [18:0] Wgt_1_752, // sfix19_En18 
  input [18:0] Wgt_1_753, // sfix19_En18 
  input [18:0] Wgt_1_754, // sfix19_En18 
  input [18:0] Wgt_1_755, // sfix19_En18 
  input [18:0] Wgt_1_756, // sfix19_En18 
  input [18:0] Wgt_1_757, // sfix19_En18 
  input [18:0] Wgt_1_758, // sfix19_En18 
  input [18:0] Wgt_1_759, // sfix19_En18 
  input [18:0] Wgt_1_760, // sfix19_En18 
  input [18:0] Wgt_1_761, // sfix19_En18 
  input [18:0] Wgt_1_762, // sfix19_En18 
  input [18:0] Wgt_1_763, // sfix19_En18 
  input [18:0] Wgt_1_764, // sfix19_En18 
  input [18:0] Wgt_1_765, // sfix19_En18 
  input [18:0] Wgt_1_766, // sfix19_En18 
  input [18:0] Wgt_1_767, // sfix19_En18 
  input [18:0] Wgt_1_768, // sfix19_En18 
  input [18:0] Wgt_1_769, // sfix19_En18 
  input [18:0] Wgt_1_770, // sfix19_En18 
  input [18:0] Wgt_1_771, // sfix19_En18 
  input [18:0] Wgt_1_772, // sfix19_En18 
  input [18:0] Wgt_1_773, // sfix19_En18 
  input [18:0] Wgt_1_774, // sfix19_En18 
  input [18:0] Wgt_1_775, // sfix19_En18 
  input [18:0] Wgt_1_776, // sfix19_En18 
  input [18:0] Wgt_1_777, // sfix19_En18 
  input [18:0] Wgt_1_778, // sfix19_En18 
  input [18:0] Wgt_1_779, // sfix19_En18 
  input [18:0] Wgt_1_780, // sfix19_En18 
  input [18:0] Wgt_1_781, // sfix19_En18 
  input [18:0] Wgt_1_782, // sfix19_En18 
  input [18:0] Wgt_1_783, // sfix19_En18 
  input [18:0] Wgt_1_784, // sfix19_En18 
  input [18:0] Wgt_2_0, // sfix19_En18 
  input [18:0] Wgt_2_1, // sfix19_En18 
  input [18:0] Wgt_2_2, // sfix19_En18 
  input [18:0] Wgt_2_3, // sfix19_En18 
  input [18:0] Wgt_2_4, // sfix19_En18 
  input [18:0] Wgt_2_5, // sfix19_En18 
  input [18:0] Wgt_2_6, // sfix19_En18 
  input [18:0] Wgt_2_7, // sfix19_En18 
  input [18:0] Wgt_2_8, // sfix19_En18 
  input [18:0] Wgt_2_9, // sfix19_En18 
  input [18:0] Wgt_2_10, // sfix19_En18 
  input [18:0] Wgt_2_11, // sfix19_En18 
  input [18:0] Wgt_2_12, // sfix19_En18 
  input [18:0] Wgt_2_13, // sfix19_En18 
  input [18:0] Wgt_2_14, // sfix19_En18 
  input [18:0] Wgt_2_15, // sfix19_En18 
  input [18:0] Wgt_2_16, // sfix19_En18 
  input [18:0] Wgt_2_17, // sfix19_En18 
  input [18:0] Wgt_2_18, // sfix19_En18 
  input [18:0] Wgt_2_19, // sfix19_En18 
  input [18:0] Wgt_2_20, // sfix19_En18 
  input [18:0] Wgt_2_21, // sfix19_En18 
  input [18:0] Wgt_2_22, // sfix19_En18 
  input [18:0] Wgt_2_23, // sfix19_En18 
  input [18:0] Wgt_2_24, // sfix19_En18 
  input [18:0] Wgt_2_25, // sfix19_En18 
  input [18:0] Wgt_2_26, // sfix19_En18 
  input [18:0] Wgt_2_27, // sfix19_En18 
  input [18:0] Wgt_2_28, // sfix19_En18 
  input [18:0] Wgt_2_29, // sfix19_En18 
  input [18:0] Wgt_2_30, // sfix19_En18 
  input [18:0] Wgt_2_31, // sfix19_En18 
  input [18:0] Wgt_2_32, // sfix19_En18 
  input [18:0] Wgt_2_33, // sfix19_En18 
  input [18:0] Wgt_2_34, // sfix19_En18 
  input [18:0] Wgt_2_35, // sfix19_En18 
  input [18:0] Wgt_2_36, // sfix19_En18 
  input [18:0] Wgt_2_37, // sfix19_En18 
  input [18:0] Wgt_2_38, // sfix19_En18 
  input [18:0] Wgt_2_39, // sfix19_En18 
  input [18:0] Wgt_2_40, // sfix19_En18 
  input [18:0] Wgt_2_41, // sfix19_En18 
  input [18:0] Wgt_2_42, // sfix19_En18 
  input [18:0] Wgt_2_43, // sfix19_En18 
  input [18:0] Wgt_2_44, // sfix19_En18 
  input [18:0] Wgt_2_45, // sfix19_En18 
  input [18:0] Wgt_2_46, // sfix19_En18 
  input [18:0] Wgt_2_47, // sfix19_En18 
  input [18:0] Wgt_2_48, // sfix19_En18 
  input [18:0] Wgt_2_49, // sfix19_En18 
  input [18:0] Wgt_2_50, // sfix19_En18 
  input [18:0] Wgt_2_51, // sfix19_En18 
  input [18:0] Wgt_2_52, // sfix19_En18 
  input [18:0] Wgt_2_53, // sfix19_En18 
  input [18:0] Wgt_2_54, // sfix19_En18 
  input [18:0] Wgt_2_55, // sfix19_En18 
  input [18:0] Wgt_2_56, // sfix19_En18 
  input [18:0] Wgt_2_57, // sfix19_En18 
  input [18:0] Wgt_2_58, // sfix19_En18 
  input [18:0] Wgt_2_59, // sfix19_En18 
  input [18:0] Wgt_2_60, // sfix19_En18 
  input [18:0] Wgt_2_61, // sfix19_En18 
  input [18:0] Wgt_2_62, // sfix19_En18 
  input [18:0] Wgt_2_63, // sfix19_En18 
  input [18:0] Wgt_2_64, // sfix19_En18 
  input [18:0] Wgt_2_65, // sfix19_En18 
  input [18:0] Wgt_2_66, // sfix19_En18 
  input [18:0] Wgt_2_67, // sfix19_En18 
  input [18:0] Wgt_2_68, // sfix19_En18 
  input [18:0] Wgt_2_69, // sfix19_En18 
  input [18:0] Wgt_2_70, // sfix19_En18 
  input [18:0] Wgt_2_71, // sfix19_En18 
  input [18:0] Wgt_2_72, // sfix19_En18 
  input [18:0] Wgt_2_73, // sfix19_En18 
  input [18:0] Wgt_2_74, // sfix19_En18 
  input [18:0] Wgt_2_75, // sfix19_En18 
  input [18:0] Wgt_2_76, // sfix19_En18 
  input [18:0] Wgt_2_77, // sfix19_En18 
  input [18:0] Wgt_2_78, // sfix19_En18 
  input [18:0] Wgt_2_79, // sfix19_En18 
  input [18:0] Wgt_2_80, // sfix19_En18 
  input [18:0] Wgt_2_81, // sfix19_En18 
  input [18:0] Wgt_2_82, // sfix19_En18 
  input [18:0] Wgt_2_83, // sfix19_En18 
  input [18:0] Wgt_2_84, // sfix19_En18 
  input [18:0] Wgt_2_85, // sfix19_En18 
  input [18:0] Wgt_2_86, // sfix19_En18 
  input [18:0] Wgt_2_87, // sfix19_En18 
  input [18:0] Wgt_2_88, // sfix19_En18 
  input [18:0] Wgt_2_89, // sfix19_En18 
  input [18:0] Wgt_2_90, // sfix19_En18 
  input [18:0] Wgt_2_91, // sfix19_En18 
  input [18:0] Wgt_2_92, // sfix19_En18 
  input [18:0] Wgt_2_93, // sfix19_En18 
  input [18:0] Wgt_2_94, // sfix19_En18 
  input [18:0] Wgt_2_95, // sfix19_En18 
  input [18:0] Wgt_2_96, // sfix19_En18 
  input [18:0] Wgt_2_97, // sfix19_En18 
  input [18:0] Wgt_2_98, // sfix19_En18 
  input [18:0] Wgt_2_99, // sfix19_En18 
  input [18:0] Wgt_2_100, // sfix19_En18 
  input [18:0] Wgt_2_101, // sfix19_En18 
  input [18:0] Wgt_2_102, // sfix19_En18 
  input [18:0] Wgt_2_103, // sfix19_En18 
  input [18:0] Wgt_2_104, // sfix19_En18 
  input [18:0] Wgt_2_105, // sfix19_En18 
  input [18:0] Wgt_2_106, // sfix19_En18 
  input [18:0] Wgt_2_107, // sfix19_En18 
  input [18:0] Wgt_2_108, // sfix19_En18 
  input [18:0] Wgt_2_109, // sfix19_En18 
  input [18:0] Wgt_2_110, // sfix19_En18 
  input [18:0] Wgt_2_111, // sfix19_En18 
  input [18:0] Wgt_2_112, // sfix19_En18 
  input [18:0] Wgt_2_113, // sfix19_En18 
  input [18:0] Wgt_2_114, // sfix19_En18 
  input [18:0] Wgt_2_115, // sfix19_En18 
  input [18:0] Wgt_2_116, // sfix19_En18 
  input [18:0] Wgt_2_117, // sfix19_En18 
  input [18:0] Wgt_2_118, // sfix19_En18 
  input [18:0] Wgt_2_119, // sfix19_En18 
  input [18:0] Wgt_2_120, // sfix19_En18 
  input [18:0] Wgt_2_121, // sfix19_En18 
  input [18:0] Wgt_2_122, // sfix19_En18 
  input [18:0] Wgt_2_123, // sfix19_En18 
  input [18:0] Wgt_2_124, // sfix19_En18 
  input [18:0] Wgt_2_125, // sfix19_En18 
  input [18:0] Wgt_2_126, // sfix19_En18 
  input [18:0] Wgt_2_127, // sfix19_En18 
  input [18:0] Wgt_2_128, // sfix19_En18 
  input [18:0] Wgt_2_129, // sfix19_En18 
  input [18:0] Wgt_2_130, // sfix19_En18 
  input [18:0] Wgt_2_131, // sfix19_En18 
  input [18:0] Wgt_2_132, // sfix19_En18 
  input [18:0] Wgt_2_133, // sfix19_En18 
  input [18:0] Wgt_2_134, // sfix19_En18 
  input [18:0] Wgt_2_135, // sfix19_En18 
  input [18:0] Wgt_2_136, // sfix19_En18 
  input [18:0] Wgt_2_137, // sfix19_En18 
  input [18:0] Wgt_2_138, // sfix19_En18 
  input [18:0] Wgt_2_139, // sfix19_En18 
  input [18:0] Wgt_2_140, // sfix19_En18 
  input [18:0] Wgt_2_141, // sfix19_En18 
  input [18:0] Wgt_2_142, // sfix19_En18 
  input [18:0] Wgt_2_143, // sfix19_En18 
  input [18:0] Wgt_2_144, // sfix19_En18 
  input [18:0] Wgt_2_145, // sfix19_En18 
  input [18:0] Wgt_2_146, // sfix19_En18 
  input [18:0] Wgt_2_147, // sfix19_En18 
  input [18:0] Wgt_2_148, // sfix19_En18 
  input [18:0] Wgt_2_149, // sfix19_En18 
  input [18:0] Wgt_2_150, // sfix19_En18 
  input [18:0] Wgt_2_151, // sfix19_En18 
  input [18:0] Wgt_2_152, // sfix19_En18 
  input [18:0] Wgt_2_153, // sfix19_En18 
  input [18:0] Wgt_2_154, // sfix19_En18 
  input [18:0] Wgt_2_155, // sfix19_En18 
  input [18:0] Wgt_2_156, // sfix19_En18 
  input [18:0] Wgt_2_157, // sfix19_En18 
  input [18:0] Wgt_2_158, // sfix19_En18 
  input [18:0] Wgt_2_159, // sfix19_En18 
  input [18:0] Wgt_2_160, // sfix19_En18 
  input [18:0] Wgt_2_161, // sfix19_En18 
  input [18:0] Wgt_2_162, // sfix19_En18 
  input [18:0] Wgt_2_163, // sfix19_En18 
  input [18:0] Wgt_2_164, // sfix19_En18 
  input [18:0] Wgt_2_165, // sfix19_En18 
  input [18:0] Wgt_2_166, // sfix19_En18 
  input [18:0] Wgt_2_167, // sfix19_En18 
  input [18:0] Wgt_2_168, // sfix19_En18 
  input [18:0] Wgt_2_169, // sfix19_En18 
  input [18:0] Wgt_2_170, // sfix19_En18 
  input [18:0] Wgt_2_171, // sfix19_En18 
  input [18:0] Wgt_2_172, // sfix19_En18 
  input [18:0] Wgt_2_173, // sfix19_En18 
  input [18:0] Wgt_2_174, // sfix19_En18 
  input [18:0] Wgt_2_175, // sfix19_En18 
  input [18:0] Wgt_2_176, // sfix19_En18 
  input [18:0] Wgt_2_177, // sfix19_En18 
  input [18:0] Wgt_2_178, // sfix19_En18 
  input [18:0] Wgt_2_179, // sfix19_En18 
  input [18:0] Wgt_2_180, // sfix19_En18 
  input [18:0] Wgt_2_181, // sfix19_En18 
  input [18:0] Wgt_2_182, // sfix19_En18 
  input [18:0] Wgt_2_183, // sfix19_En18 
  input [18:0] Wgt_2_184, // sfix19_En18 
  input [18:0] Wgt_2_185, // sfix19_En18 
  input [18:0] Wgt_2_186, // sfix19_En18 
  input [18:0] Wgt_2_187, // sfix19_En18 
  input [18:0] Wgt_2_188, // sfix19_En18 
  input [18:0] Wgt_2_189, // sfix19_En18 
  input [18:0] Wgt_2_190, // sfix19_En18 
  input [18:0] Wgt_2_191, // sfix19_En18 
  input [18:0] Wgt_2_192, // sfix19_En18 
  input [18:0] Wgt_2_193, // sfix19_En18 
  input [18:0] Wgt_2_194, // sfix19_En18 
  input [18:0] Wgt_2_195, // sfix19_En18 
  input [18:0] Wgt_2_196, // sfix19_En18 
  input [18:0] Wgt_2_197, // sfix19_En18 
  input [18:0] Wgt_2_198, // sfix19_En18 
  input [18:0] Wgt_2_199, // sfix19_En18 
  input [18:0] Wgt_2_200, // sfix19_En18 
  input [18:0] Wgt_2_201, // sfix19_En18 
  input [18:0] Wgt_2_202, // sfix19_En18 
  input [18:0] Wgt_2_203, // sfix19_En18 
  input [18:0] Wgt_2_204, // sfix19_En18 
  input [18:0] Wgt_2_205, // sfix19_En18 
  input [18:0] Wgt_2_206, // sfix19_En18 
  input [18:0] Wgt_2_207, // sfix19_En18 
  input [18:0] Wgt_2_208, // sfix19_En18 
  input [18:0] Wgt_2_209, // sfix19_En18 
  input [18:0] Wgt_2_210, // sfix19_En18 
  input [18:0] Wgt_2_211, // sfix19_En18 
  input [18:0] Wgt_2_212, // sfix19_En18 
  input [18:0] Wgt_2_213, // sfix19_En18 
  input [18:0] Wgt_2_214, // sfix19_En18 
  input [18:0] Wgt_2_215, // sfix19_En18 
  input [18:0] Wgt_2_216, // sfix19_En18 
  input [18:0] Wgt_2_217, // sfix19_En18 
  input [18:0] Wgt_2_218, // sfix19_En18 
  input [18:0] Wgt_2_219, // sfix19_En18 
  input [18:0] Wgt_2_220, // sfix19_En18 
  input [18:0] Wgt_2_221, // sfix19_En18 
  input [18:0] Wgt_2_222, // sfix19_En18 
  input [18:0] Wgt_2_223, // sfix19_En18 
  input [18:0] Wgt_2_224, // sfix19_En18 
  input [18:0] Wgt_2_225, // sfix19_En18 
  input [18:0] Wgt_2_226, // sfix19_En18 
  input [18:0] Wgt_2_227, // sfix19_En18 
  input [18:0] Wgt_2_228, // sfix19_En18 
  input [18:0] Wgt_2_229, // sfix19_En18 
  input [18:0] Wgt_2_230, // sfix19_En18 
  input [18:0] Wgt_2_231, // sfix19_En18 
  input [18:0] Wgt_2_232, // sfix19_En18 
  input [18:0] Wgt_2_233, // sfix19_En18 
  input [18:0] Wgt_2_234, // sfix19_En18 
  input [18:0] Wgt_2_235, // sfix19_En18 
  input [18:0] Wgt_2_236, // sfix19_En18 
  input [18:0] Wgt_2_237, // sfix19_En18 
  input [18:0] Wgt_2_238, // sfix19_En18 
  input [18:0] Wgt_2_239, // sfix19_En18 
  input [18:0] Wgt_2_240, // sfix19_En18 
  input [18:0] Wgt_2_241, // sfix19_En18 
  input [18:0] Wgt_2_242, // sfix19_En18 
  input [18:0] Wgt_2_243, // sfix19_En18 
  input [18:0] Wgt_2_244, // sfix19_En18 
  input [18:0] Wgt_2_245, // sfix19_En18 
  input [18:0] Wgt_2_246, // sfix19_En18 
  input [18:0] Wgt_2_247, // sfix19_En18 
  input [18:0] Wgt_2_248, // sfix19_En18 
  input [18:0] Wgt_2_249, // sfix19_En18 
  input [18:0] Wgt_2_250, // sfix19_En18 
  input [18:0] Wgt_2_251, // sfix19_En18 
  input [18:0] Wgt_2_252, // sfix19_En18 
  input [18:0] Wgt_2_253, // sfix19_En18 
  input [18:0] Wgt_2_254, // sfix19_En18 
  input [18:0] Wgt_2_255, // sfix19_En18 
  input [18:0] Wgt_2_256, // sfix19_En18 
  input [18:0] Wgt_2_257, // sfix19_En18 
  input [18:0] Wgt_2_258, // sfix19_En18 
  input [18:0] Wgt_2_259, // sfix19_En18 
  input [18:0] Wgt_2_260, // sfix19_En18 
  input [18:0] Wgt_2_261, // sfix19_En18 
  input [18:0] Wgt_2_262, // sfix19_En18 
  input [18:0] Wgt_2_263, // sfix19_En18 
  input [18:0] Wgt_2_264, // sfix19_En18 
  input [18:0] Wgt_2_265, // sfix19_En18 
  input [18:0] Wgt_2_266, // sfix19_En18 
  input [18:0] Wgt_2_267, // sfix19_En18 
  input [18:0] Wgt_2_268, // sfix19_En18 
  input [18:0] Wgt_2_269, // sfix19_En18 
  input [18:0] Wgt_2_270, // sfix19_En18 
  input [18:0] Wgt_2_271, // sfix19_En18 
  input [18:0] Wgt_2_272, // sfix19_En18 
  input [18:0] Wgt_2_273, // sfix19_En18 
  input [18:0] Wgt_2_274, // sfix19_En18 
  input [18:0] Wgt_2_275, // sfix19_En18 
  input [18:0] Wgt_2_276, // sfix19_En18 
  input [18:0] Wgt_2_277, // sfix19_En18 
  input [18:0] Wgt_2_278, // sfix19_En18 
  input [18:0] Wgt_2_279, // sfix19_En18 
  input [18:0] Wgt_2_280, // sfix19_En18 
  input [18:0] Wgt_2_281, // sfix19_En18 
  input [18:0] Wgt_2_282, // sfix19_En18 
  input [18:0] Wgt_2_283, // sfix19_En18 
  input [18:0] Wgt_2_284, // sfix19_En18 
  input [18:0] Wgt_2_285, // sfix19_En18 
  input [18:0] Wgt_2_286, // sfix19_En18 
  input [18:0] Wgt_2_287, // sfix19_En18 
  input [18:0] Wgt_2_288, // sfix19_En18 
  input [18:0] Wgt_2_289, // sfix19_En18 
  input [18:0] Wgt_2_290, // sfix19_En18 
  input [18:0] Wgt_2_291, // sfix19_En18 
  input [18:0] Wgt_2_292, // sfix19_En18 
  input [18:0] Wgt_2_293, // sfix19_En18 
  input [18:0] Wgt_2_294, // sfix19_En18 
  input [18:0] Wgt_2_295, // sfix19_En18 
  input [18:0] Wgt_2_296, // sfix19_En18 
  input [18:0] Wgt_2_297, // sfix19_En18 
  input [18:0] Wgt_2_298, // sfix19_En18 
  input [18:0] Wgt_2_299, // sfix19_En18 
  input [18:0] Wgt_2_300, // sfix19_En18 
  input [18:0] Wgt_2_301, // sfix19_En18 
  input [18:0] Wgt_2_302, // sfix19_En18 
  input [18:0] Wgt_2_303, // sfix19_En18 
  input [18:0] Wgt_2_304, // sfix19_En18 
  input [18:0] Wgt_2_305, // sfix19_En18 
  input [18:0] Wgt_2_306, // sfix19_En18 
  input [18:0] Wgt_2_307, // sfix19_En18 
  input [18:0] Wgt_2_308, // sfix19_En18 
  input [18:0] Wgt_2_309, // sfix19_En18 
  input [18:0] Wgt_2_310, // sfix19_En18 
  input [18:0] Wgt_2_311, // sfix19_En18 
  input [18:0] Wgt_2_312, // sfix19_En18 
  input [18:0] Wgt_2_313, // sfix19_En18 
  input [18:0] Wgt_2_314, // sfix19_En18 
  input [18:0] Wgt_2_315, // sfix19_En18 
  input [18:0] Wgt_2_316, // sfix19_En18 
  input [18:0] Wgt_2_317, // sfix19_En18 
  input [18:0] Wgt_2_318, // sfix19_En18 
  input [18:0] Wgt_2_319, // sfix19_En18 
  input [18:0] Wgt_2_320, // sfix19_En18 
  input [18:0] Wgt_2_321, // sfix19_En18 
  input [18:0] Wgt_2_322, // sfix19_En18 
  input [18:0] Wgt_2_323, // sfix19_En18 
  input [18:0] Wgt_2_324, // sfix19_En18 
  input [18:0] Wgt_2_325, // sfix19_En18 
  input [18:0] Wgt_2_326, // sfix19_En18 
  input [18:0] Wgt_2_327, // sfix19_En18 
  input [18:0] Wgt_2_328, // sfix19_En18 
  input [18:0] Wgt_2_329, // sfix19_En18 
  input [18:0] Wgt_2_330, // sfix19_En18 
  input [18:0] Wgt_2_331, // sfix19_En18 
  input [18:0] Wgt_2_332, // sfix19_En18 
  input [18:0] Wgt_2_333, // sfix19_En18 
  input [18:0] Wgt_2_334, // sfix19_En18 
  input [18:0] Wgt_2_335, // sfix19_En18 
  input [18:0] Wgt_2_336, // sfix19_En18 
  input [18:0] Wgt_2_337, // sfix19_En18 
  input [18:0] Wgt_2_338, // sfix19_En18 
  input [18:0] Wgt_2_339, // sfix19_En18 
  input [18:0] Wgt_2_340, // sfix19_En18 
  input [18:0] Wgt_2_341, // sfix19_En18 
  input [18:0] Wgt_2_342, // sfix19_En18 
  input [18:0] Wgt_2_343, // sfix19_En18 
  input [18:0] Wgt_2_344, // sfix19_En18 
  input [18:0] Wgt_2_345, // sfix19_En18 
  input [18:0] Wgt_2_346, // sfix19_En18 
  input [18:0] Wgt_2_347, // sfix19_En18 
  input [18:0] Wgt_2_348, // sfix19_En18 
  input [18:0] Wgt_2_349, // sfix19_En18 
  input [18:0] Wgt_2_350, // sfix19_En18 
  input [18:0] Wgt_2_351, // sfix19_En18 
  input [18:0] Wgt_2_352, // sfix19_En18 
  input [18:0] Wgt_2_353, // sfix19_En18 
  input [18:0] Wgt_2_354, // sfix19_En18 
  input [18:0] Wgt_2_355, // sfix19_En18 
  input [18:0] Wgt_2_356, // sfix19_En18 
  input [18:0] Wgt_2_357, // sfix19_En18 
  input [18:0] Wgt_2_358, // sfix19_En18 
  input [18:0] Wgt_2_359, // sfix19_En18 
  input [18:0] Wgt_2_360, // sfix19_En18 
  input [18:0] Wgt_2_361, // sfix19_En18 
  input [18:0] Wgt_2_362, // sfix19_En18 
  input [18:0] Wgt_2_363, // sfix19_En18 
  input [18:0] Wgt_2_364, // sfix19_En18 
  input [18:0] Wgt_2_365, // sfix19_En18 
  input [18:0] Wgt_2_366, // sfix19_En18 
  input [18:0] Wgt_2_367, // sfix19_En18 
  input [18:0] Wgt_2_368, // sfix19_En18 
  input [18:0] Wgt_2_369, // sfix19_En18 
  input [18:0] Wgt_2_370, // sfix19_En18 
  input [18:0] Wgt_2_371, // sfix19_En18 
  input [18:0] Wgt_2_372, // sfix19_En18 
  input [18:0] Wgt_2_373, // sfix19_En18 
  input [18:0] Wgt_2_374, // sfix19_En18 
  input [18:0] Wgt_2_375, // sfix19_En18 
  input [18:0] Wgt_2_376, // sfix19_En18 
  input [18:0] Wgt_2_377, // sfix19_En18 
  input [18:0] Wgt_2_378, // sfix19_En18 
  input [18:0] Wgt_2_379, // sfix19_En18 
  input [18:0] Wgt_2_380, // sfix19_En18 
  input [18:0] Wgt_2_381, // sfix19_En18 
  input [18:0] Wgt_2_382, // sfix19_En18 
  input [18:0] Wgt_2_383, // sfix19_En18 
  input [18:0] Wgt_2_384, // sfix19_En18 
  input [18:0] Wgt_2_385, // sfix19_En18 
  input [18:0] Wgt_2_386, // sfix19_En18 
  input [18:0] Wgt_2_387, // sfix19_En18 
  input [18:0] Wgt_2_388, // sfix19_En18 
  input [18:0] Wgt_2_389, // sfix19_En18 
  input [18:0] Wgt_2_390, // sfix19_En18 
  input [18:0] Wgt_2_391, // sfix19_En18 
  input [18:0] Wgt_2_392, // sfix19_En18 
  input [18:0] Wgt_2_393, // sfix19_En18 
  input [18:0] Wgt_2_394, // sfix19_En18 
  input [18:0] Wgt_2_395, // sfix19_En18 
  input [18:0] Wgt_2_396, // sfix19_En18 
  input [18:0] Wgt_2_397, // sfix19_En18 
  input [18:0] Wgt_2_398, // sfix19_En18 
  input [18:0] Wgt_2_399, // sfix19_En18 
  input [18:0] Wgt_2_400, // sfix19_En18 
  input [18:0] Wgt_2_401, // sfix19_En18 
  input [18:0] Wgt_2_402, // sfix19_En18 
  input [18:0] Wgt_2_403, // sfix19_En18 
  input [18:0] Wgt_2_404, // sfix19_En18 
  input [18:0] Wgt_2_405, // sfix19_En18 
  input [18:0] Wgt_2_406, // sfix19_En18 
  input [18:0] Wgt_2_407, // sfix19_En18 
  input [18:0] Wgt_2_408, // sfix19_En18 
  input [18:0] Wgt_2_409, // sfix19_En18 
  input [18:0] Wgt_2_410, // sfix19_En18 
  input [18:0] Wgt_2_411, // sfix19_En18 
  input [18:0] Wgt_2_412, // sfix19_En18 
  input [18:0] Wgt_2_413, // sfix19_En18 
  input [18:0] Wgt_2_414, // sfix19_En18 
  input [18:0] Wgt_2_415, // sfix19_En18 
  input [18:0] Wgt_2_416, // sfix19_En18 
  input [18:0] Wgt_2_417, // sfix19_En18 
  input [18:0] Wgt_2_418, // sfix19_En18 
  input [18:0] Wgt_2_419, // sfix19_En18 
  input [18:0] Wgt_2_420, // sfix19_En18 
  input [18:0] Wgt_2_421, // sfix19_En18 
  input [18:0] Wgt_2_422, // sfix19_En18 
  input [18:0] Wgt_2_423, // sfix19_En18 
  input [18:0] Wgt_2_424, // sfix19_En18 
  input [18:0] Wgt_2_425, // sfix19_En18 
  input [18:0] Wgt_2_426, // sfix19_En18 
  input [18:0] Wgt_2_427, // sfix19_En18 
  input [18:0] Wgt_2_428, // sfix19_En18 
  input [18:0] Wgt_2_429, // sfix19_En18 
  input [18:0] Wgt_2_430, // sfix19_En18 
  input [18:0] Wgt_2_431, // sfix19_En18 
  input [18:0] Wgt_2_432, // sfix19_En18 
  input [18:0] Wgt_2_433, // sfix19_En18 
  input [18:0] Wgt_2_434, // sfix19_En18 
  input [18:0] Wgt_2_435, // sfix19_En18 
  input [18:0] Wgt_2_436, // sfix19_En18 
  input [18:0] Wgt_2_437, // sfix19_En18 
  input [18:0] Wgt_2_438, // sfix19_En18 
  input [18:0] Wgt_2_439, // sfix19_En18 
  input [18:0] Wgt_2_440, // sfix19_En18 
  input [18:0] Wgt_2_441, // sfix19_En18 
  input [18:0] Wgt_2_442, // sfix19_En18 
  input [18:0] Wgt_2_443, // sfix19_En18 
  input [18:0] Wgt_2_444, // sfix19_En18 
  input [18:0] Wgt_2_445, // sfix19_En18 
  input [18:0] Wgt_2_446, // sfix19_En18 
  input [18:0] Wgt_2_447, // sfix19_En18 
  input [18:0] Wgt_2_448, // sfix19_En18 
  input [18:0] Wgt_2_449, // sfix19_En18 
  input [18:0] Wgt_2_450, // sfix19_En18 
  input [18:0] Wgt_2_451, // sfix19_En18 
  input [18:0] Wgt_2_452, // sfix19_En18 
  input [18:0] Wgt_2_453, // sfix19_En18 
  input [18:0] Wgt_2_454, // sfix19_En18 
  input [18:0] Wgt_2_455, // sfix19_En18 
  input [18:0] Wgt_2_456, // sfix19_En18 
  input [18:0] Wgt_2_457, // sfix19_En18 
  input [18:0] Wgt_2_458, // sfix19_En18 
  input [18:0] Wgt_2_459, // sfix19_En18 
  input [18:0] Wgt_2_460, // sfix19_En18 
  input [18:0] Wgt_2_461, // sfix19_En18 
  input [18:0] Wgt_2_462, // sfix19_En18 
  input [18:0] Wgt_2_463, // sfix19_En18 
  input [18:0] Wgt_2_464, // sfix19_En18 
  input [18:0] Wgt_2_465, // sfix19_En18 
  input [18:0] Wgt_2_466, // sfix19_En18 
  input [18:0] Wgt_2_467, // sfix19_En18 
  input [18:0] Wgt_2_468, // sfix19_En18 
  input [18:0] Wgt_2_469, // sfix19_En18 
  input [18:0] Wgt_2_470, // sfix19_En18 
  input [18:0] Wgt_2_471, // sfix19_En18 
  input [18:0] Wgt_2_472, // sfix19_En18 
  input [18:0] Wgt_2_473, // sfix19_En18 
  input [18:0] Wgt_2_474, // sfix19_En18 
  input [18:0] Wgt_2_475, // sfix19_En18 
  input [18:0] Wgt_2_476, // sfix19_En18 
  input [18:0] Wgt_2_477, // sfix19_En18 
  input [18:0] Wgt_2_478, // sfix19_En18 
  input [18:0] Wgt_2_479, // sfix19_En18 
  input [18:0] Wgt_2_480, // sfix19_En18 
  input [18:0] Wgt_2_481, // sfix19_En18 
  input [18:0] Wgt_2_482, // sfix19_En18 
  input [18:0] Wgt_2_483, // sfix19_En18 
  input [18:0] Wgt_2_484, // sfix19_En18 
  input [18:0] Wgt_2_485, // sfix19_En18 
  input [18:0] Wgt_2_486, // sfix19_En18 
  input [18:0] Wgt_2_487, // sfix19_En18 
  input [18:0] Wgt_2_488, // sfix19_En18 
  input [18:0] Wgt_2_489, // sfix19_En18 
  input [18:0] Wgt_2_490, // sfix19_En18 
  input [18:0] Wgt_2_491, // sfix19_En18 
  input [18:0] Wgt_2_492, // sfix19_En18 
  input [18:0] Wgt_2_493, // sfix19_En18 
  input [18:0] Wgt_2_494, // sfix19_En18 
  input [18:0] Wgt_2_495, // sfix19_En18 
  input [18:0] Wgt_2_496, // sfix19_En18 
  input [18:0] Wgt_2_497, // sfix19_En18 
  input [18:0] Wgt_2_498, // sfix19_En18 
  input [18:0] Wgt_2_499, // sfix19_En18 
  input [18:0] Wgt_2_500, // sfix19_En18 
  input [18:0] Wgt_2_501, // sfix19_En18 
  input [18:0] Wgt_2_502, // sfix19_En18 
  input [18:0] Wgt_2_503, // sfix19_En18 
  input [18:0] Wgt_2_504, // sfix19_En18 
  input [18:0] Wgt_2_505, // sfix19_En18 
  input [18:0] Wgt_2_506, // sfix19_En18 
  input [18:0] Wgt_2_507, // sfix19_En18 
  input [18:0] Wgt_2_508, // sfix19_En18 
  input [18:0] Wgt_2_509, // sfix19_En18 
  input [18:0] Wgt_2_510, // sfix19_En18 
  input [18:0] Wgt_2_511, // sfix19_En18 
  input [18:0] Wgt_2_512, // sfix19_En18 
  input [18:0] Wgt_2_513, // sfix19_En18 
  input [18:0] Wgt_2_514, // sfix19_En18 
  input [18:0] Wgt_2_515, // sfix19_En18 
  input [18:0] Wgt_2_516, // sfix19_En18 
  input [18:0] Wgt_2_517, // sfix19_En18 
  input [18:0] Wgt_2_518, // sfix19_En18 
  input [18:0] Wgt_2_519, // sfix19_En18 
  input [18:0] Wgt_2_520, // sfix19_En18 
  input [18:0] Wgt_2_521, // sfix19_En18 
  input [18:0] Wgt_2_522, // sfix19_En18 
  input [18:0] Wgt_2_523, // sfix19_En18 
  input [18:0] Wgt_2_524, // sfix19_En18 
  input [18:0] Wgt_2_525, // sfix19_En18 
  input [18:0] Wgt_2_526, // sfix19_En18 
  input [18:0] Wgt_2_527, // sfix19_En18 
  input [18:0] Wgt_2_528, // sfix19_En18 
  input [18:0] Wgt_2_529, // sfix19_En18 
  input [18:0] Wgt_2_530, // sfix19_En18 
  input [18:0] Wgt_2_531, // sfix19_En18 
  input [18:0] Wgt_2_532, // sfix19_En18 
  input [18:0] Wgt_2_533, // sfix19_En18 
  input [18:0] Wgt_2_534, // sfix19_En18 
  input [18:0] Wgt_2_535, // sfix19_En18 
  input [18:0] Wgt_2_536, // sfix19_En18 
  input [18:0] Wgt_2_537, // sfix19_En18 
  input [18:0] Wgt_2_538, // sfix19_En18 
  input [18:0] Wgt_2_539, // sfix19_En18 
  input [18:0] Wgt_2_540, // sfix19_En18 
  input [18:0] Wgt_2_541, // sfix19_En18 
  input [18:0] Wgt_2_542, // sfix19_En18 
  input [18:0] Wgt_2_543, // sfix19_En18 
  input [18:0] Wgt_2_544, // sfix19_En18 
  input [18:0] Wgt_2_545, // sfix19_En18 
  input [18:0] Wgt_2_546, // sfix19_En18 
  input [18:0] Wgt_2_547, // sfix19_En18 
  input [18:0] Wgt_2_548, // sfix19_En18 
  input [18:0] Wgt_2_549, // sfix19_En18 
  input [18:0] Wgt_2_550, // sfix19_En18 
  input [18:0] Wgt_2_551, // sfix19_En18 
  input [18:0] Wgt_2_552, // sfix19_En18 
  input [18:0] Wgt_2_553, // sfix19_En18 
  input [18:0] Wgt_2_554, // sfix19_En18 
  input [18:0] Wgt_2_555, // sfix19_En18 
  input [18:0] Wgt_2_556, // sfix19_En18 
  input [18:0] Wgt_2_557, // sfix19_En18 
  input [18:0] Wgt_2_558, // sfix19_En18 
  input [18:0] Wgt_2_559, // sfix19_En18 
  input [18:0] Wgt_2_560, // sfix19_En18 
  input [18:0] Wgt_2_561, // sfix19_En18 
  input [18:0] Wgt_2_562, // sfix19_En18 
  input [18:0] Wgt_2_563, // sfix19_En18 
  input [18:0] Wgt_2_564, // sfix19_En18 
  input [18:0] Wgt_2_565, // sfix19_En18 
  input [18:0] Wgt_2_566, // sfix19_En18 
  input [18:0] Wgt_2_567, // sfix19_En18 
  input [18:0] Wgt_2_568, // sfix19_En18 
  input [18:0] Wgt_2_569, // sfix19_En18 
  input [18:0] Wgt_2_570, // sfix19_En18 
  input [18:0] Wgt_2_571, // sfix19_En18 
  input [18:0] Wgt_2_572, // sfix19_En18 
  input [18:0] Wgt_2_573, // sfix19_En18 
  input [18:0] Wgt_2_574, // sfix19_En18 
  input [18:0] Wgt_2_575, // sfix19_En18 
  input [18:0] Wgt_2_576, // sfix19_En18 
  input [18:0] Wgt_2_577, // sfix19_En18 
  input [18:0] Wgt_2_578, // sfix19_En18 
  input [18:0] Wgt_2_579, // sfix19_En18 
  input [18:0] Wgt_2_580, // sfix19_En18 
  input [18:0] Wgt_2_581, // sfix19_En18 
  input [18:0] Wgt_2_582, // sfix19_En18 
  input [18:0] Wgt_2_583, // sfix19_En18 
  input [18:0] Wgt_2_584, // sfix19_En18 
  input [18:0] Wgt_2_585, // sfix19_En18 
  input [18:0] Wgt_2_586, // sfix19_En18 
  input [18:0] Wgt_2_587, // sfix19_En18 
  input [18:0] Wgt_2_588, // sfix19_En18 
  input [18:0] Wgt_2_589, // sfix19_En18 
  input [18:0] Wgt_2_590, // sfix19_En18 
  input [18:0] Wgt_2_591, // sfix19_En18 
  input [18:0] Wgt_2_592, // sfix19_En18 
  input [18:0] Wgt_2_593, // sfix19_En18 
  input [18:0] Wgt_2_594, // sfix19_En18 
  input [18:0] Wgt_2_595, // sfix19_En18 
  input [18:0] Wgt_2_596, // sfix19_En18 
  input [18:0] Wgt_2_597, // sfix19_En18 
  input [18:0] Wgt_2_598, // sfix19_En18 
  input [18:0] Wgt_2_599, // sfix19_En18 
  input [18:0] Wgt_2_600, // sfix19_En18 
  input [18:0] Wgt_2_601, // sfix19_En18 
  input [18:0] Wgt_2_602, // sfix19_En18 
  input [18:0] Wgt_2_603, // sfix19_En18 
  input [18:0] Wgt_2_604, // sfix19_En18 
  input [18:0] Wgt_2_605, // sfix19_En18 
  input [18:0] Wgt_2_606, // sfix19_En18 
  input [18:0] Wgt_2_607, // sfix19_En18 
  input [18:0] Wgt_2_608, // sfix19_En18 
  input [18:0] Wgt_2_609, // sfix19_En18 
  input [18:0] Wgt_2_610, // sfix19_En18 
  input [18:0] Wgt_2_611, // sfix19_En18 
  input [18:0] Wgt_2_612, // sfix19_En18 
  input [18:0] Wgt_2_613, // sfix19_En18 
  input [18:0] Wgt_2_614, // sfix19_En18 
  input [18:0] Wgt_2_615, // sfix19_En18 
  input [18:0] Wgt_2_616, // sfix19_En18 
  input [18:0] Wgt_2_617, // sfix19_En18 
  input [18:0] Wgt_2_618, // sfix19_En18 
  input [18:0] Wgt_2_619, // sfix19_En18 
  input [18:0] Wgt_2_620, // sfix19_En18 
  input [18:0] Wgt_2_621, // sfix19_En18 
  input [18:0] Wgt_2_622, // sfix19_En18 
  input [18:0] Wgt_2_623, // sfix19_En18 
  input [18:0] Wgt_2_624, // sfix19_En18 
  input [18:0] Wgt_2_625, // sfix19_En18 
  input [18:0] Wgt_2_626, // sfix19_En18 
  input [18:0] Wgt_2_627, // sfix19_En18 
  input [18:0] Wgt_2_628, // sfix19_En18 
  input [18:0] Wgt_2_629, // sfix19_En18 
  input [18:0] Wgt_2_630, // sfix19_En18 
  input [18:0] Wgt_2_631, // sfix19_En18 
  input [18:0] Wgt_2_632, // sfix19_En18 
  input [18:0] Wgt_2_633, // sfix19_En18 
  input [18:0] Wgt_2_634, // sfix19_En18 
  input [18:0] Wgt_2_635, // sfix19_En18 
  input [18:0] Wgt_2_636, // sfix19_En18 
  input [18:0] Wgt_2_637, // sfix19_En18 
  input [18:0] Wgt_2_638, // sfix19_En18 
  input [18:0] Wgt_2_639, // sfix19_En18 
  input [18:0] Wgt_2_640, // sfix19_En18 
  input [18:0] Wgt_2_641, // sfix19_En18 
  input [18:0] Wgt_2_642, // sfix19_En18 
  input [18:0] Wgt_2_643, // sfix19_En18 
  input [18:0] Wgt_2_644, // sfix19_En18 
  input [18:0] Wgt_2_645, // sfix19_En18 
  input [18:0] Wgt_2_646, // sfix19_En18 
  input [18:0] Wgt_2_647, // sfix19_En18 
  input [18:0] Wgt_2_648, // sfix19_En18 
  input [18:0] Wgt_2_649, // sfix19_En18 
  input [18:0] Wgt_2_650, // sfix19_En18 
  input [18:0] Wgt_2_651, // sfix19_En18 
  input [18:0] Wgt_2_652, // sfix19_En18 
  input [18:0] Wgt_2_653, // sfix19_En18 
  input [18:0] Wgt_2_654, // sfix19_En18 
  input [18:0] Wgt_2_655, // sfix19_En18 
  input [18:0] Wgt_2_656, // sfix19_En18 
  input [18:0] Wgt_2_657, // sfix19_En18 
  input [18:0] Wgt_2_658, // sfix19_En18 
  input [18:0] Wgt_2_659, // sfix19_En18 
  input [18:0] Wgt_2_660, // sfix19_En18 
  input [18:0] Wgt_2_661, // sfix19_En18 
  input [18:0] Wgt_2_662, // sfix19_En18 
  input [18:0] Wgt_2_663, // sfix19_En18 
  input [18:0] Wgt_2_664, // sfix19_En18 
  input [18:0] Wgt_2_665, // sfix19_En18 
  input [18:0] Wgt_2_666, // sfix19_En18 
  input [18:0] Wgt_2_667, // sfix19_En18 
  input [18:0] Wgt_2_668, // sfix19_En18 
  input [18:0] Wgt_2_669, // sfix19_En18 
  input [18:0] Wgt_2_670, // sfix19_En18 
  input [18:0] Wgt_2_671, // sfix19_En18 
  input [18:0] Wgt_2_672, // sfix19_En18 
  input [18:0] Wgt_2_673, // sfix19_En18 
  input [18:0] Wgt_2_674, // sfix19_En18 
  input [18:0] Wgt_2_675, // sfix19_En18 
  input [18:0] Wgt_2_676, // sfix19_En18 
  input [18:0] Wgt_2_677, // sfix19_En18 
  input [18:0] Wgt_2_678, // sfix19_En18 
  input [18:0] Wgt_2_679, // sfix19_En18 
  input [18:0] Wgt_2_680, // sfix19_En18 
  input [18:0] Wgt_2_681, // sfix19_En18 
  input [18:0] Wgt_2_682, // sfix19_En18 
  input [18:0] Wgt_2_683, // sfix19_En18 
  input [18:0] Wgt_2_684, // sfix19_En18 
  input [18:0] Wgt_2_685, // sfix19_En18 
  input [18:0] Wgt_2_686, // sfix19_En18 
  input [18:0] Wgt_2_687, // sfix19_En18 
  input [18:0] Wgt_2_688, // sfix19_En18 
  input [18:0] Wgt_2_689, // sfix19_En18 
  input [18:0] Wgt_2_690, // sfix19_En18 
  input [18:0] Wgt_2_691, // sfix19_En18 
  input [18:0] Wgt_2_692, // sfix19_En18 
  input [18:0] Wgt_2_693, // sfix19_En18 
  input [18:0] Wgt_2_694, // sfix19_En18 
  input [18:0] Wgt_2_695, // sfix19_En18 
  input [18:0] Wgt_2_696, // sfix19_En18 
  input [18:0] Wgt_2_697, // sfix19_En18 
  input [18:0] Wgt_2_698, // sfix19_En18 
  input [18:0] Wgt_2_699, // sfix19_En18 
  input [18:0] Wgt_2_700, // sfix19_En18 
  input [18:0] Wgt_2_701, // sfix19_En18 
  input [18:0] Wgt_2_702, // sfix19_En18 
  input [18:0] Wgt_2_703, // sfix19_En18 
  input [18:0] Wgt_2_704, // sfix19_En18 
  input [18:0] Wgt_2_705, // sfix19_En18 
  input [18:0] Wgt_2_706, // sfix19_En18 
  input [18:0] Wgt_2_707, // sfix19_En18 
  input [18:0] Wgt_2_708, // sfix19_En18 
  input [18:0] Wgt_2_709, // sfix19_En18 
  input [18:0] Wgt_2_710, // sfix19_En18 
  input [18:0] Wgt_2_711, // sfix19_En18 
  input [18:0] Wgt_2_712, // sfix19_En18 
  input [18:0] Wgt_2_713, // sfix19_En18 
  input [18:0] Wgt_2_714, // sfix19_En18 
  input [18:0] Wgt_2_715, // sfix19_En18 
  input [18:0] Wgt_2_716, // sfix19_En18 
  input [18:0] Wgt_2_717, // sfix19_En18 
  input [18:0] Wgt_2_718, // sfix19_En18 
  input [18:0] Wgt_2_719, // sfix19_En18 
  input [18:0] Wgt_2_720, // sfix19_En18 
  input [18:0] Wgt_2_721, // sfix19_En18 
  input [18:0] Wgt_2_722, // sfix19_En18 
  input [18:0] Wgt_2_723, // sfix19_En18 
  input [18:0] Wgt_2_724, // sfix19_En18 
  input [18:0] Wgt_2_725, // sfix19_En18 
  input [18:0] Wgt_2_726, // sfix19_En18 
  input [18:0] Wgt_2_727, // sfix19_En18 
  input [18:0] Wgt_2_728, // sfix19_En18 
  input [18:0] Wgt_2_729, // sfix19_En18 
  input [18:0] Wgt_2_730, // sfix19_En18 
  input [18:0] Wgt_2_731, // sfix19_En18 
  input [18:0] Wgt_2_732, // sfix19_En18 
  input [18:0] Wgt_2_733, // sfix19_En18 
  input [18:0] Wgt_2_734, // sfix19_En18 
  input [18:0] Wgt_2_735, // sfix19_En18 
  input [18:0] Wgt_2_736, // sfix19_En18 
  input [18:0] Wgt_2_737, // sfix19_En18 
  input [18:0] Wgt_2_738, // sfix19_En18 
  input [18:0] Wgt_2_739, // sfix19_En18 
  input [18:0] Wgt_2_740, // sfix19_En18 
  input [18:0] Wgt_2_741, // sfix19_En18 
  input [18:0] Wgt_2_742, // sfix19_En18 
  input [18:0] Wgt_2_743, // sfix19_En18 
  input [18:0] Wgt_2_744, // sfix19_En18 
  input [18:0] Wgt_2_745, // sfix19_En18 
  input [18:0] Wgt_2_746, // sfix19_En18 
  input [18:0] Wgt_2_747, // sfix19_En18 
  input [18:0] Wgt_2_748, // sfix19_En18 
  input [18:0] Wgt_2_749, // sfix19_En18 
  input [18:0] Wgt_2_750, // sfix19_En18 
  input [18:0] Wgt_2_751, // sfix19_En18 
  input [18:0] Wgt_2_752, // sfix19_En18 
  input [18:0] Wgt_2_753, // sfix19_En18 
  input [18:0] Wgt_2_754, // sfix19_En18 
  input [18:0] Wgt_2_755, // sfix19_En18 
  input [18:0] Wgt_2_756, // sfix19_En18 
  input [18:0] Wgt_2_757, // sfix19_En18 
  input [18:0] Wgt_2_758, // sfix19_En18 
  input [18:0] Wgt_2_759, // sfix19_En18 
  input [18:0] Wgt_2_760, // sfix19_En18 
  input [18:0] Wgt_2_761, // sfix19_En18 
  input [18:0] Wgt_2_762, // sfix19_En18 
  input [18:0] Wgt_2_763, // sfix19_En18 
  input [18:0] Wgt_2_764, // sfix19_En18 
  input [18:0] Wgt_2_765, // sfix19_En18 
  input [18:0] Wgt_2_766, // sfix19_En18 
  input [18:0] Wgt_2_767, // sfix19_En18 
  input [18:0] Wgt_2_768, // sfix19_En18 
  input [18:0] Wgt_2_769, // sfix19_En18 
  input [18:0] Wgt_2_770, // sfix19_En18 
  input [18:0] Wgt_2_771, // sfix19_En18 
  input [18:0] Wgt_2_772, // sfix19_En18 
  input [18:0] Wgt_2_773, // sfix19_En18 
  input [18:0] Wgt_2_774, // sfix19_En18 
  input [18:0] Wgt_2_775, // sfix19_En18 
  input [18:0] Wgt_2_776, // sfix19_En18 
  input [18:0] Wgt_2_777, // sfix19_En18 
  input [18:0] Wgt_2_778, // sfix19_En18 
  input [18:0] Wgt_2_779, // sfix19_En18 
  input [18:0] Wgt_2_780, // sfix19_En18 
  input [18:0] Wgt_2_781, // sfix19_En18 
  input [18:0] Wgt_2_782, // sfix19_En18 
  input [18:0] Wgt_2_783, // sfix19_En18 
  input [18:0] Wgt_2_784, // sfix19_En18 
  input [18:0] Wgt_3_0, // sfix19_En18 
  input [18:0] Wgt_3_1, // sfix19_En18 
  input [18:0] Wgt_3_2, // sfix19_En18 
  input [18:0] Wgt_3_3, // sfix19_En18 
  input [18:0] Wgt_3_4, // sfix19_En18 
  input [18:0] Wgt_3_5, // sfix19_En18 
  input [18:0] Wgt_3_6, // sfix19_En18 
  input [18:0] Wgt_3_7, // sfix19_En18 
  input [18:0] Wgt_3_8, // sfix19_En18 
  input [18:0] Wgt_3_9, // sfix19_En18 
  input [18:0] Wgt_3_10, // sfix19_En18 
  input [18:0] Wgt_3_11, // sfix19_En18 
  input [18:0] Wgt_3_12, // sfix19_En18 
  input [18:0] Wgt_3_13, // sfix19_En18 
  input [18:0] Wgt_3_14, // sfix19_En18 
  input [18:0] Wgt_3_15, // sfix19_En18 
  input [18:0] Wgt_3_16, // sfix19_En18 
  input [18:0] Wgt_3_17, // sfix19_En18 
  input [18:0] Wgt_3_18, // sfix19_En18 
  input [18:0] Wgt_3_19, // sfix19_En18 
  input [18:0] Wgt_3_20, // sfix19_En18 
  input [18:0] Wgt_3_21, // sfix19_En18 
  input [18:0] Wgt_3_22, // sfix19_En18 
  input [18:0] Wgt_3_23, // sfix19_En18 
  input [18:0] Wgt_3_24, // sfix19_En18 
  input [18:0] Wgt_3_25, // sfix19_En18 
  input [18:0] Wgt_3_26, // sfix19_En18 
  input [18:0] Wgt_3_27, // sfix19_En18 
  input [18:0] Wgt_3_28, // sfix19_En18 
  input [18:0] Wgt_3_29, // sfix19_En18 
  input [18:0] Wgt_3_30, // sfix19_En18 
  input [18:0] Wgt_3_31, // sfix19_En18 
  input [18:0] Wgt_3_32, // sfix19_En18 
  input [18:0] Wgt_3_33, // sfix19_En18 
  input [18:0] Wgt_3_34, // sfix19_En18 
  input [18:0] Wgt_3_35, // sfix19_En18 
  input [18:0] Wgt_3_36, // sfix19_En18 
  input [18:0] Wgt_3_37, // sfix19_En18 
  input [18:0] Wgt_3_38, // sfix19_En18 
  input [18:0] Wgt_3_39, // sfix19_En18 
  input [18:0] Wgt_3_40, // sfix19_En18 
  input [18:0] Wgt_3_41, // sfix19_En18 
  input [18:0] Wgt_3_42, // sfix19_En18 
  input [18:0] Wgt_3_43, // sfix19_En18 
  input [18:0] Wgt_3_44, // sfix19_En18 
  input [18:0] Wgt_3_45, // sfix19_En18 
  input [18:0] Wgt_3_46, // sfix19_En18 
  input [18:0] Wgt_3_47, // sfix19_En18 
  input [18:0] Wgt_3_48, // sfix19_En18 
  input [18:0] Wgt_3_49, // sfix19_En18 
  input [18:0] Wgt_3_50, // sfix19_En18 
  input [18:0] Wgt_3_51, // sfix19_En18 
  input [18:0] Wgt_3_52, // sfix19_En18 
  input [18:0] Wgt_3_53, // sfix19_En18 
  input [18:0] Wgt_3_54, // sfix19_En18 
  input [18:0] Wgt_3_55, // sfix19_En18 
  input [18:0] Wgt_3_56, // sfix19_En18 
  input [18:0] Wgt_3_57, // sfix19_En18 
  input [18:0] Wgt_3_58, // sfix19_En18 
  input [18:0] Wgt_3_59, // sfix19_En18 
  input [18:0] Wgt_3_60, // sfix19_En18 
  input [18:0] Wgt_3_61, // sfix19_En18 
  input [18:0] Wgt_3_62, // sfix19_En18 
  input [18:0] Wgt_3_63, // sfix19_En18 
  input [18:0] Wgt_3_64, // sfix19_En18 
  input [18:0] Wgt_3_65, // sfix19_En18 
  input [18:0] Wgt_3_66, // sfix19_En18 
  input [18:0] Wgt_3_67, // sfix19_En18 
  input [18:0] Wgt_3_68, // sfix19_En18 
  input [18:0] Wgt_3_69, // sfix19_En18 
  input [18:0] Wgt_3_70, // sfix19_En18 
  input [18:0] Wgt_3_71, // sfix19_En18 
  input [18:0] Wgt_3_72, // sfix19_En18 
  input [18:0] Wgt_3_73, // sfix19_En18 
  input [18:0] Wgt_3_74, // sfix19_En18 
  input [18:0] Wgt_3_75, // sfix19_En18 
  input [18:0] Wgt_3_76, // sfix19_En18 
  input [18:0] Wgt_3_77, // sfix19_En18 
  input [18:0] Wgt_3_78, // sfix19_En18 
  input [18:0] Wgt_3_79, // sfix19_En18 
  input [18:0] Wgt_3_80, // sfix19_En18 
  input [18:0] Wgt_3_81, // sfix19_En18 
  input [18:0] Wgt_3_82, // sfix19_En18 
  input [18:0] Wgt_3_83, // sfix19_En18 
  input [18:0] Wgt_3_84, // sfix19_En18 
  input [18:0] Wgt_3_85, // sfix19_En18 
  input [18:0] Wgt_3_86, // sfix19_En18 
  input [18:0] Wgt_3_87, // sfix19_En18 
  input [18:0] Wgt_3_88, // sfix19_En18 
  input [18:0] Wgt_3_89, // sfix19_En18 
  input [18:0] Wgt_3_90, // sfix19_En18 
  input [18:0] Wgt_3_91, // sfix19_En18 
  input [18:0] Wgt_3_92, // sfix19_En18 
  input [18:0] Wgt_3_93, // sfix19_En18 
  input [18:0] Wgt_3_94, // sfix19_En18 
  input [18:0] Wgt_3_95, // sfix19_En18 
  input [18:0] Wgt_3_96, // sfix19_En18 
  input [18:0] Wgt_3_97, // sfix19_En18 
  input [18:0] Wgt_3_98, // sfix19_En18 
  input [18:0] Wgt_3_99, // sfix19_En18 
  input [18:0] Wgt_3_100, // sfix19_En18 
  input [18:0] Wgt_3_101, // sfix19_En18 
  input [18:0] Wgt_3_102, // sfix19_En18 
  input [18:0] Wgt_3_103, // sfix19_En18 
  input [18:0] Wgt_3_104, // sfix19_En18 
  input [18:0] Wgt_3_105, // sfix19_En18 
  input [18:0] Wgt_3_106, // sfix19_En18 
  input [18:0] Wgt_3_107, // sfix19_En18 
  input [18:0] Wgt_3_108, // sfix19_En18 
  input [18:0] Wgt_3_109, // sfix19_En18 
  input [18:0] Wgt_3_110, // sfix19_En18 
  input [18:0] Wgt_3_111, // sfix19_En18 
  input [18:0] Wgt_3_112, // sfix19_En18 
  input [18:0] Wgt_3_113, // sfix19_En18 
  input [18:0] Wgt_3_114, // sfix19_En18 
  input [18:0] Wgt_3_115, // sfix19_En18 
  input [18:0] Wgt_3_116, // sfix19_En18 
  input [18:0] Wgt_3_117, // sfix19_En18 
  input [18:0] Wgt_3_118, // sfix19_En18 
  input [18:0] Wgt_3_119, // sfix19_En18 
  input [18:0] Wgt_3_120, // sfix19_En18 
  input [18:0] Wgt_3_121, // sfix19_En18 
  input [18:0] Wgt_3_122, // sfix19_En18 
  input [18:0] Wgt_3_123, // sfix19_En18 
  input [18:0] Wgt_3_124, // sfix19_En18 
  input [18:0] Wgt_3_125, // sfix19_En18 
  input [18:0] Wgt_3_126, // sfix19_En18 
  input [18:0] Wgt_3_127, // sfix19_En18 
  input [18:0] Wgt_3_128, // sfix19_En18 
  input [18:0] Wgt_3_129, // sfix19_En18 
  input [18:0] Wgt_3_130, // sfix19_En18 
  input [18:0] Wgt_3_131, // sfix19_En18 
  input [18:0] Wgt_3_132, // sfix19_En18 
  input [18:0] Wgt_3_133, // sfix19_En18 
  input [18:0] Wgt_3_134, // sfix19_En18 
  input [18:0] Wgt_3_135, // sfix19_En18 
  input [18:0] Wgt_3_136, // sfix19_En18 
  input [18:0] Wgt_3_137, // sfix19_En18 
  input [18:0] Wgt_3_138, // sfix19_En18 
  input [18:0] Wgt_3_139, // sfix19_En18 
  input [18:0] Wgt_3_140, // sfix19_En18 
  input [18:0] Wgt_3_141, // sfix19_En18 
  input [18:0] Wgt_3_142, // sfix19_En18 
  input [18:0] Wgt_3_143, // sfix19_En18 
  input [18:0] Wgt_3_144, // sfix19_En18 
  input [18:0] Wgt_3_145, // sfix19_En18 
  input [18:0] Wgt_3_146, // sfix19_En18 
  input [18:0] Wgt_3_147, // sfix19_En18 
  input [18:0] Wgt_3_148, // sfix19_En18 
  input [18:0] Wgt_3_149, // sfix19_En18 
  input [18:0] Wgt_3_150, // sfix19_En18 
  input [18:0] Wgt_3_151, // sfix19_En18 
  input [18:0] Wgt_3_152, // sfix19_En18 
  input [18:0] Wgt_3_153, // sfix19_En18 
  input [18:0] Wgt_3_154, // sfix19_En18 
  input [18:0] Wgt_3_155, // sfix19_En18 
  input [18:0] Wgt_3_156, // sfix19_En18 
  input [18:0] Wgt_3_157, // sfix19_En18 
  input [18:0] Wgt_3_158, // sfix19_En18 
  input [18:0] Wgt_3_159, // sfix19_En18 
  input [18:0] Wgt_3_160, // sfix19_En18 
  input [18:0] Wgt_3_161, // sfix19_En18 
  input [18:0] Wgt_3_162, // sfix19_En18 
  input [18:0] Wgt_3_163, // sfix19_En18 
  input [18:0] Wgt_3_164, // sfix19_En18 
  input [18:0] Wgt_3_165, // sfix19_En18 
  input [18:0] Wgt_3_166, // sfix19_En18 
  input [18:0] Wgt_3_167, // sfix19_En18 
  input [18:0] Wgt_3_168, // sfix19_En18 
  input [18:0] Wgt_3_169, // sfix19_En18 
  input [18:0] Wgt_3_170, // sfix19_En18 
  input [18:0] Wgt_3_171, // sfix19_En18 
  input [18:0] Wgt_3_172, // sfix19_En18 
  input [18:0] Wgt_3_173, // sfix19_En18 
  input [18:0] Wgt_3_174, // sfix19_En18 
  input [18:0] Wgt_3_175, // sfix19_En18 
  input [18:0] Wgt_3_176, // sfix19_En18 
  input [18:0] Wgt_3_177, // sfix19_En18 
  input [18:0] Wgt_3_178, // sfix19_En18 
  input [18:0] Wgt_3_179, // sfix19_En18 
  input [18:0] Wgt_3_180, // sfix19_En18 
  input [18:0] Wgt_3_181, // sfix19_En18 
  input [18:0] Wgt_3_182, // sfix19_En18 
  input [18:0] Wgt_3_183, // sfix19_En18 
  input [18:0] Wgt_3_184, // sfix19_En18 
  input [18:0] Wgt_3_185, // sfix19_En18 
  input [18:0] Wgt_3_186, // sfix19_En18 
  input [18:0] Wgt_3_187, // sfix19_En18 
  input [18:0] Wgt_3_188, // sfix19_En18 
  input [18:0] Wgt_3_189, // sfix19_En18 
  input [18:0] Wgt_3_190, // sfix19_En18 
  input [18:0] Wgt_3_191, // sfix19_En18 
  input [18:0] Wgt_3_192, // sfix19_En18 
  input [18:0] Wgt_3_193, // sfix19_En18 
  input [18:0] Wgt_3_194, // sfix19_En18 
  input [18:0] Wgt_3_195, // sfix19_En18 
  input [18:0] Wgt_3_196, // sfix19_En18 
  input [18:0] Wgt_3_197, // sfix19_En18 
  input [18:0] Wgt_3_198, // sfix19_En18 
  input [18:0] Wgt_3_199, // sfix19_En18 
  input [18:0] Wgt_3_200, // sfix19_En18 
  input [18:0] Wgt_3_201, // sfix19_En18 
  input [18:0] Wgt_3_202, // sfix19_En18 
  input [18:0] Wgt_3_203, // sfix19_En18 
  input [18:0] Wgt_3_204, // sfix19_En18 
  input [18:0] Wgt_3_205, // sfix19_En18 
  input [18:0] Wgt_3_206, // sfix19_En18 
  input [18:0] Wgt_3_207, // sfix19_En18 
  input [18:0] Wgt_3_208, // sfix19_En18 
  input [18:0] Wgt_3_209, // sfix19_En18 
  input [18:0] Wgt_3_210, // sfix19_En18 
  input [18:0] Wgt_3_211, // sfix19_En18 
  input [18:0] Wgt_3_212, // sfix19_En18 
  input [18:0] Wgt_3_213, // sfix19_En18 
  input [18:0] Wgt_3_214, // sfix19_En18 
  input [18:0] Wgt_3_215, // sfix19_En18 
  input [18:0] Wgt_3_216, // sfix19_En18 
  input [18:0] Wgt_3_217, // sfix19_En18 
  input [18:0] Wgt_3_218, // sfix19_En18 
  input [18:0] Wgt_3_219, // sfix19_En18 
  input [18:0] Wgt_3_220, // sfix19_En18 
  input [18:0] Wgt_3_221, // sfix19_En18 
  input [18:0] Wgt_3_222, // sfix19_En18 
  input [18:0] Wgt_3_223, // sfix19_En18 
  input [18:0] Wgt_3_224, // sfix19_En18 
  input [18:0] Wgt_3_225, // sfix19_En18 
  input [18:0] Wgt_3_226, // sfix19_En18 
  input [18:0] Wgt_3_227, // sfix19_En18 
  input [18:0] Wgt_3_228, // sfix19_En18 
  input [18:0] Wgt_3_229, // sfix19_En18 
  input [18:0] Wgt_3_230, // sfix19_En18 
  input [18:0] Wgt_3_231, // sfix19_En18 
  input [18:0] Wgt_3_232, // sfix19_En18 
  input [18:0] Wgt_3_233, // sfix19_En18 
  input [18:0] Wgt_3_234, // sfix19_En18 
  input [18:0] Wgt_3_235, // sfix19_En18 
  input [18:0] Wgt_3_236, // sfix19_En18 
  input [18:0] Wgt_3_237, // sfix19_En18 
  input [18:0] Wgt_3_238, // sfix19_En18 
  input [18:0] Wgt_3_239, // sfix19_En18 
  input [18:0] Wgt_3_240, // sfix19_En18 
  input [18:0] Wgt_3_241, // sfix19_En18 
  input [18:0] Wgt_3_242, // sfix19_En18 
  input [18:0] Wgt_3_243, // sfix19_En18 
  input [18:0] Wgt_3_244, // sfix19_En18 
  input [18:0] Wgt_3_245, // sfix19_En18 
  input [18:0] Wgt_3_246, // sfix19_En18 
  input [18:0] Wgt_3_247, // sfix19_En18 
  input [18:0] Wgt_3_248, // sfix19_En18 
  input [18:0] Wgt_3_249, // sfix19_En18 
  input [18:0] Wgt_3_250, // sfix19_En18 
  input [18:0] Wgt_3_251, // sfix19_En18 
  input [18:0] Wgt_3_252, // sfix19_En18 
  input [18:0] Wgt_3_253, // sfix19_En18 
  input [18:0] Wgt_3_254, // sfix19_En18 
  input [18:0] Wgt_3_255, // sfix19_En18 
  input [18:0] Wgt_3_256, // sfix19_En18 
  input [18:0] Wgt_3_257, // sfix19_En18 
  input [18:0] Wgt_3_258, // sfix19_En18 
  input [18:0] Wgt_3_259, // sfix19_En18 
  input [18:0] Wgt_3_260, // sfix19_En18 
  input [18:0] Wgt_3_261, // sfix19_En18 
  input [18:0] Wgt_3_262, // sfix19_En18 
  input [18:0] Wgt_3_263, // sfix19_En18 
  input [18:0] Wgt_3_264, // sfix19_En18 
  input [18:0] Wgt_3_265, // sfix19_En18 
  input [18:0] Wgt_3_266, // sfix19_En18 
  input [18:0] Wgt_3_267, // sfix19_En18 
  input [18:0] Wgt_3_268, // sfix19_En18 
  input [18:0] Wgt_3_269, // sfix19_En18 
  input [18:0] Wgt_3_270, // sfix19_En18 
  input [18:0] Wgt_3_271, // sfix19_En18 
  input [18:0] Wgt_3_272, // sfix19_En18 
  input [18:0] Wgt_3_273, // sfix19_En18 
  input [18:0] Wgt_3_274, // sfix19_En18 
  input [18:0] Wgt_3_275, // sfix19_En18 
  input [18:0] Wgt_3_276, // sfix19_En18 
  input [18:0] Wgt_3_277, // sfix19_En18 
  input [18:0] Wgt_3_278, // sfix19_En18 
  input [18:0] Wgt_3_279, // sfix19_En18 
  input [18:0] Wgt_3_280, // sfix19_En18 
  input [18:0] Wgt_3_281, // sfix19_En18 
  input [18:0] Wgt_3_282, // sfix19_En18 
  input [18:0] Wgt_3_283, // sfix19_En18 
  input [18:0] Wgt_3_284, // sfix19_En18 
  input [18:0] Wgt_3_285, // sfix19_En18 
  input [18:0] Wgt_3_286, // sfix19_En18 
  input [18:0] Wgt_3_287, // sfix19_En18 
  input [18:0] Wgt_3_288, // sfix19_En18 
  input [18:0] Wgt_3_289, // sfix19_En18 
  input [18:0] Wgt_3_290, // sfix19_En18 
  input [18:0] Wgt_3_291, // sfix19_En18 
  input [18:0] Wgt_3_292, // sfix19_En18 
  input [18:0] Wgt_3_293, // sfix19_En18 
  input [18:0] Wgt_3_294, // sfix19_En18 
  input [18:0] Wgt_3_295, // sfix19_En18 
  input [18:0] Wgt_3_296, // sfix19_En18 
  input [18:0] Wgt_3_297, // sfix19_En18 
  input [18:0] Wgt_3_298, // sfix19_En18 
  input [18:0] Wgt_3_299, // sfix19_En18 
  input [18:0] Wgt_3_300, // sfix19_En18 
  input [18:0] Wgt_3_301, // sfix19_En18 
  input [18:0] Wgt_3_302, // sfix19_En18 
  input [18:0] Wgt_3_303, // sfix19_En18 
  input [18:0] Wgt_3_304, // sfix19_En18 
  input [18:0] Wgt_3_305, // sfix19_En18 
  input [18:0] Wgt_3_306, // sfix19_En18 
  input [18:0] Wgt_3_307, // sfix19_En18 
  input [18:0] Wgt_3_308, // sfix19_En18 
  input [18:0] Wgt_3_309, // sfix19_En18 
  input [18:0] Wgt_3_310, // sfix19_En18 
  input [18:0] Wgt_3_311, // sfix19_En18 
  input [18:0] Wgt_3_312, // sfix19_En18 
  input [18:0] Wgt_3_313, // sfix19_En18 
  input [18:0] Wgt_3_314, // sfix19_En18 
  input [18:0] Wgt_3_315, // sfix19_En18 
  input [18:0] Wgt_3_316, // sfix19_En18 
  input [18:0] Wgt_3_317, // sfix19_En18 
  input [18:0] Wgt_3_318, // sfix19_En18 
  input [18:0] Wgt_3_319, // sfix19_En18 
  input [18:0] Wgt_3_320, // sfix19_En18 
  input [18:0] Wgt_3_321, // sfix19_En18 
  input [18:0] Wgt_3_322, // sfix19_En18 
  input [18:0] Wgt_3_323, // sfix19_En18 
  input [18:0] Wgt_3_324, // sfix19_En18 
  input [18:0] Wgt_3_325, // sfix19_En18 
  input [18:0] Wgt_3_326, // sfix19_En18 
  input [18:0] Wgt_3_327, // sfix19_En18 
  input [18:0] Wgt_3_328, // sfix19_En18 
  input [18:0] Wgt_3_329, // sfix19_En18 
  input [18:0] Wgt_3_330, // sfix19_En18 
  input [18:0] Wgt_3_331, // sfix19_En18 
  input [18:0] Wgt_3_332, // sfix19_En18 
  input [18:0] Wgt_3_333, // sfix19_En18 
  input [18:0] Wgt_3_334, // sfix19_En18 
  input [18:0] Wgt_3_335, // sfix19_En18 
  input [18:0] Wgt_3_336, // sfix19_En18 
  input [18:0] Wgt_3_337, // sfix19_En18 
  input [18:0] Wgt_3_338, // sfix19_En18 
  input [18:0] Wgt_3_339, // sfix19_En18 
  input [18:0] Wgt_3_340, // sfix19_En18 
  input [18:0] Wgt_3_341, // sfix19_En18 
  input [18:0] Wgt_3_342, // sfix19_En18 
  input [18:0] Wgt_3_343, // sfix19_En18 
  input [18:0] Wgt_3_344, // sfix19_En18 
  input [18:0] Wgt_3_345, // sfix19_En18 
  input [18:0] Wgt_3_346, // sfix19_En18 
  input [18:0] Wgt_3_347, // sfix19_En18 
  input [18:0] Wgt_3_348, // sfix19_En18 
  input [18:0] Wgt_3_349, // sfix19_En18 
  input [18:0] Wgt_3_350, // sfix19_En18 
  input [18:0] Wgt_3_351, // sfix19_En18 
  input [18:0] Wgt_3_352, // sfix19_En18 
  input [18:0] Wgt_3_353, // sfix19_En18 
  input [18:0] Wgt_3_354, // sfix19_En18 
  input [18:0] Wgt_3_355, // sfix19_En18 
  input [18:0] Wgt_3_356, // sfix19_En18 
  input [18:0] Wgt_3_357, // sfix19_En18 
  input [18:0] Wgt_3_358, // sfix19_En18 
  input [18:0] Wgt_3_359, // sfix19_En18 
  input [18:0] Wgt_3_360, // sfix19_En18 
  input [18:0] Wgt_3_361, // sfix19_En18 
  input [18:0] Wgt_3_362, // sfix19_En18 
  input [18:0] Wgt_3_363, // sfix19_En18 
  input [18:0] Wgt_3_364, // sfix19_En18 
  input [18:0] Wgt_3_365, // sfix19_En18 
  input [18:0] Wgt_3_366, // sfix19_En18 
  input [18:0] Wgt_3_367, // sfix19_En18 
  input [18:0] Wgt_3_368, // sfix19_En18 
  input [18:0] Wgt_3_369, // sfix19_En18 
  input [18:0] Wgt_3_370, // sfix19_En18 
  input [18:0] Wgt_3_371, // sfix19_En18 
  input [18:0] Wgt_3_372, // sfix19_En18 
  input [18:0] Wgt_3_373, // sfix19_En18 
  input [18:0] Wgt_3_374, // sfix19_En18 
  input [18:0] Wgt_3_375, // sfix19_En18 
  input [18:0] Wgt_3_376, // sfix19_En18 
  input [18:0] Wgt_3_377, // sfix19_En18 
  input [18:0] Wgt_3_378, // sfix19_En18 
  input [18:0] Wgt_3_379, // sfix19_En18 
  input [18:0] Wgt_3_380, // sfix19_En18 
  input [18:0] Wgt_3_381, // sfix19_En18 
  input [18:0] Wgt_3_382, // sfix19_En18 
  input [18:0] Wgt_3_383, // sfix19_En18 
  input [18:0] Wgt_3_384, // sfix19_En18 
  input [18:0] Wgt_3_385, // sfix19_En18 
  input [18:0] Wgt_3_386, // sfix19_En18 
  input [18:0] Wgt_3_387, // sfix19_En18 
  input [18:0] Wgt_3_388, // sfix19_En18 
  input [18:0] Wgt_3_389, // sfix19_En18 
  input [18:0] Wgt_3_390, // sfix19_En18 
  input [18:0] Wgt_3_391, // sfix19_En18 
  input [18:0] Wgt_3_392, // sfix19_En18 
  input [18:0] Wgt_3_393, // sfix19_En18 
  input [18:0] Wgt_3_394, // sfix19_En18 
  input [18:0] Wgt_3_395, // sfix19_En18 
  input [18:0] Wgt_3_396, // sfix19_En18 
  input [18:0] Wgt_3_397, // sfix19_En18 
  input [18:0] Wgt_3_398, // sfix19_En18 
  input [18:0] Wgt_3_399, // sfix19_En18 
  input [18:0] Wgt_3_400, // sfix19_En18 
  input [18:0] Wgt_3_401, // sfix19_En18 
  input [18:0] Wgt_3_402, // sfix19_En18 
  input [18:0] Wgt_3_403, // sfix19_En18 
  input [18:0] Wgt_3_404, // sfix19_En18 
  input [18:0] Wgt_3_405, // sfix19_En18 
  input [18:0] Wgt_3_406, // sfix19_En18 
  input [18:0] Wgt_3_407, // sfix19_En18 
  input [18:0] Wgt_3_408, // sfix19_En18 
  input [18:0] Wgt_3_409, // sfix19_En18 
  input [18:0] Wgt_3_410, // sfix19_En18 
  input [18:0] Wgt_3_411, // sfix19_En18 
  input [18:0] Wgt_3_412, // sfix19_En18 
  input [18:0] Wgt_3_413, // sfix19_En18 
  input [18:0] Wgt_3_414, // sfix19_En18 
  input [18:0] Wgt_3_415, // sfix19_En18 
  input [18:0] Wgt_3_416, // sfix19_En18 
  input [18:0] Wgt_3_417, // sfix19_En18 
  input [18:0] Wgt_3_418, // sfix19_En18 
  input [18:0] Wgt_3_419, // sfix19_En18 
  input [18:0] Wgt_3_420, // sfix19_En18 
  input [18:0] Wgt_3_421, // sfix19_En18 
  input [18:0] Wgt_3_422, // sfix19_En18 
  input [18:0] Wgt_3_423, // sfix19_En18 
  input [18:0] Wgt_3_424, // sfix19_En18 
  input [18:0] Wgt_3_425, // sfix19_En18 
  input [18:0] Wgt_3_426, // sfix19_En18 
  input [18:0] Wgt_3_427, // sfix19_En18 
  input [18:0] Wgt_3_428, // sfix19_En18 
  input [18:0] Wgt_3_429, // sfix19_En18 
  input [18:0] Wgt_3_430, // sfix19_En18 
  input [18:0] Wgt_3_431, // sfix19_En18 
  input [18:0] Wgt_3_432, // sfix19_En18 
  input [18:0] Wgt_3_433, // sfix19_En18 
  input [18:0] Wgt_3_434, // sfix19_En18 
  input [18:0] Wgt_3_435, // sfix19_En18 
  input [18:0] Wgt_3_436, // sfix19_En18 
  input [18:0] Wgt_3_437, // sfix19_En18 
  input [18:0] Wgt_3_438, // sfix19_En18 
  input [18:0] Wgt_3_439, // sfix19_En18 
  input [18:0] Wgt_3_440, // sfix19_En18 
  input [18:0] Wgt_3_441, // sfix19_En18 
  input [18:0] Wgt_3_442, // sfix19_En18 
  input [18:0] Wgt_3_443, // sfix19_En18 
  input [18:0] Wgt_3_444, // sfix19_En18 
  input [18:0] Wgt_3_445, // sfix19_En18 
  input [18:0] Wgt_3_446, // sfix19_En18 
  input [18:0] Wgt_3_447, // sfix19_En18 
  input [18:0] Wgt_3_448, // sfix19_En18 
  input [18:0] Wgt_3_449, // sfix19_En18 
  input [18:0] Wgt_3_450, // sfix19_En18 
  input [18:0] Wgt_3_451, // sfix19_En18 
  input [18:0] Wgt_3_452, // sfix19_En18 
  input [18:0] Wgt_3_453, // sfix19_En18 
  input [18:0] Wgt_3_454, // sfix19_En18 
  input [18:0] Wgt_3_455, // sfix19_En18 
  input [18:0] Wgt_3_456, // sfix19_En18 
  input [18:0] Wgt_3_457, // sfix19_En18 
  input [18:0] Wgt_3_458, // sfix19_En18 
  input [18:0] Wgt_3_459, // sfix19_En18 
  input [18:0] Wgt_3_460, // sfix19_En18 
  input [18:0] Wgt_3_461, // sfix19_En18 
  input [18:0] Wgt_3_462, // sfix19_En18 
  input [18:0] Wgt_3_463, // sfix19_En18 
  input [18:0] Wgt_3_464, // sfix19_En18 
  input [18:0] Wgt_3_465, // sfix19_En18 
  input [18:0] Wgt_3_466, // sfix19_En18 
  input [18:0] Wgt_3_467, // sfix19_En18 
  input [18:0] Wgt_3_468, // sfix19_En18 
  input [18:0] Wgt_3_469, // sfix19_En18 
  input [18:0] Wgt_3_470, // sfix19_En18 
  input [18:0] Wgt_3_471, // sfix19_En18 
  input [18:0] Wgt_3_472, // sfix19_En18 
  input [18:0] Wgt_3_473, // sfix19_En18 
  input [18:0] Wgt_3_474, // sfix19_En18 
  input [18:0] Wgt_3_475, // sfix19_En18 
  input [18:0] Wgt_3_476, // sfix19_En18 
  input [18:0] Wgt_3_477, // sfix19_En18 
  input [18:0] Wgt_3_478, // sfix19_En18 
  input [18:0] Wgt_3_479, // sfix19_En18 
  input [18:0] Wgt_3_480, // sfix19_En18 
  input [18:0] Wgt_3_481, // sfix19_En18 
  input [18:0] Wgt_3_482, // sfix19_En18 
  input [18:0] Wgt_3_483, // sfix19_En18 
  input [18:0] Wgt_3_484, // sfix19_En18 
  input [18:0] Wgt_3_485, // sfix19_En18 
  input [18:0] Wgt_3_486, // sfix19_En18 
  input [18:0] Wgt_3_487, // sfix19_En18 
  input [18:0] Wgt_3_488, // sfix19_En18 
  input [18:0] Wgt_3_489, // sfix19_En18 
  input [18:0] Wgt_3_490, // sfix19_En18 
  input [18:0] Wgt_3_491, // sfix19_En18 
  input [18:0] Wgt_3_492, // sfix19_En18 
  input [18:0] Wgt_3_493, // sfix19_En18 
  input [18:0] Wgt_3_494, // sfix19_En18 
  input [18:0] Wgt_3_495, // sfix19_En18 
  input [18:0] Wgt_3_496, // sfix19_En18 
  input [18:0] Wgt_3_497, // sfix19_En18 
  input [18:0] Wgt_3_498, // sfix19_En18 
  input [18:0] Wgt_3_499, // sfix19_En18 
  input [18:0] Wgt_3_500, // sfix19_En18 
  input [18:0] Wgt_3_501, // sfix19_En18 
  input [18:0] Wgt_3_502, // sfix19_En18 
  input [18:0] Wgt_3_503, // sfix19_En18 
  input [18:0] Wgt_3_504, // sfix19_En18 
  input [18:0] Wgt_3_505, // sfix19_En18 
  input [18:0] Wgt_3_506, // sfix19_En18 
  input [18:0] Wgt_3_507, // sfix19_En18 
  input [18:0] Wgt_3_508, // sfix19_En18 
  input [18:0] Wgt_3_509, // sfix19_En18 
  input [18:0] Wgt_3_510, // sfix19_En18 
  input [18:0] Wgt_3_511, // sfix19_En18 
  input [18:0] Wgt_3_512, // sfix19_En18 
  input [18:0] Wgt_3_513, // sfix19_En18 
  input [18:0] Wgt_3_514, // sfix19_En18 
  input [18:0] Wgt_3_515, // sfix19_En18 
  input [18:0] Wgt_3_516, // sfix19_En18 
  input [18:0] Wgt_3_517, // sfix19_En18 
  input [18:0] Wgt_3_518, // sfix19_En18 
  input [18:0] Wgt_3_519, // sfix19_En18 
  input [18:0] Wgt_3_520, // sfix19_En18 
  input [18:0] Wgt_3_521, // sfix19_En18 
  input [18:0] Wgt_3_522, // sfix19_En18 
  input [18:0] Wgt_3_523, // sfix19_En18 
  input [18:0] Wgt_3_524, // sfix19_En18 
  input [18:0] Wgt_3_525, // sfix19_En18 
  input [18:0] Wgt_3_526, // sfix19_En18 
  input [18:0] Wgt_3_527, // sfix19_En18 
  input [18:0] Wgt_3_528, // sfix19_En18 
  input [18:0] Wgt_3_529, // sfix19_En18 
  input [18:0] Wgt_3_530, // sfix19_En18 
  input [18:0] Wgt_3_531, // sfix19_En18 
  input [18:0] Wgt_3_532, // sfix19_En18 
  input [18:0] Wgt_3_533, // sfix19_En18 
  input [18:0] Wgt_3_534, // sfix19_En18 
  input [18:0] Wgt_3_535, // sfix19_En18 
  input [18:0] Wgt_3_536, // sfix19_En18 
  input [18:0] Wgt_3_537, // sfix19_En18 
  input [18:0] Wgt_3_538, // sfix19_En18 
  input [18:0] Wgt_3_539, // sfix19_En18 
  input [18:0] Wgt_3_540, // sfix19_En18 
  input [18:0] Wgt_3_541, // sfix19_En18 
  input [18:0] Wgt_3_542, // sfix19_En18 
  input [18:0] Wgt_3_543, // sfix19_En18 
  input [18:0] Wgt_3_544, // sfix19_En18 
  input [18:0] Wgt_3_545, // sfix19_En18 
  input [18:0] Wgt_3_546, // sfix19_En18 
  input [18:0] Wgt_3_547, // sfix19_En18 
  input [18:0] Wgt_3_548, // sfix19_En18 
  input [18:0] Wgt_3_549, // sfix19_En18 
  input [18:0] Wgt_3_550, // sfix19_En18 
  input [18:0] Wgt_3_551, // sfix19_En18 
  input [18:0] Wgt_3_552, // sfix19_En18 
  input [18:0] Wgt_3_553, // sfix19_En18 
  input [18:0] Wgt_3_554, // sfix19_En18 
  input [18:0] Wgt_3_555, // sfix19_En18 
  input [18:0] Wgt_3_556, // sfix19_En18 
  input [18:0] Wgt_3_557, // sfix19_En18 
  input [18:0] Wgt_3_558, // sfix19_En18 
  input [18:0] Wgt_3_559, // sfix19_En18 
  input [18:0] Wgt_3_560, // sfix19_En18 
  input [18:0] Wgt_3_561, // sfix19_En18 
  input [18:0] Wgt_3_562, // sfix19_En18 
  input [18:0] Wgt_3_563, // sfix19_En18 
  input [18:0] Wgt_3_564, // sfix19_En18 
  input [18:0] Wgt_3_565, // sfix19_En18 
  input [18:0] Wgt_3_566, // sfix19_En18 
  input [18:0] Wgt_3_567, // sfix19_En18 
  input [18:0] Wgt_3_568, // sfix19_En18 
  input [18:0] Wgt_3_569, // sfix19_En18 
  input [18:0] Wgt_3_570, // sfix19_En18 
  input [18:0] Wgt_3_571, // sfix19_En18 
  input [18:0] Wgt_3_572, // sfix19_En18 
  input [18:0] Wgt_3_573, // sfix19_En18 
  input [18:0] Wgt_3_574, // sfix19_En18 
  input [18:0] Wgt_3_575, // sfix19_En18 
  input [18:0] Wgt_3_576, // sfix19_En18 
  input [18:0] Wgt_3_577, // sfix19_En18 
  input [18:0] Wgt_3_578, // sfix19_En18 
  input [18:0] Wgt_3_579, // sfix19_En18 
  input [18:0] Wgt_3_580, // sfix19_En18 
  input [18:0] Wgt_3_581, // sfix19_En18 
  input [18:0] Wgt_3_582, // sfix19_En18 
  input [18:0] Wgt_3_583, // sfix19_En18 
  input [18:0] Wgt_3_584, // sfix19_En18 
  input [18:0] Wgt_3_585, // sfix19_En18 
  input [18:0] Wgt_3_586, // sfix19_En18 
  input [18:0] Wgt_3_587, // sfix19_En18 
  input [18:0] Wgt_3_588, // sfix19_En18 
  input [18:0] Wgt_3_589, // sfix19_En18 
  input [18:0] Wgt_3_590, // sfix19_En18 
  input [18:0] Wgt_3_591, // sfix19_En18 
  input [18:0] Wgt_3_592, // sfix19_En18 
  input [18:0] Wgt_3_593, // sfix19_En18 
  input [18:0] Wgt_3_594, // sfix19_En18 
  input [18:0] Wgt_3_595, // sfix19_En18 
  input [18:0] Wgt_3_596, // sfix19_En18 
  input [18:0] Wgt_3_597, // sfix19_En18 
  input [18:0] Wgt_3_598, // sfix19_En18 
  input [18:0] Wgt_3_599, // sfix19_En18 
  input [18:0] Wgt_3_600, // sfix19_En18 
  input [18:0] Wgt_3_601, // sfix19_En18 
  input [18:0] Wgt_3_602, // sfix19_En18 
  input [18:0] Wgt_3_603, // sfix19_En18 
  input [18:0] Wgt_3_604, // sfix19_En18 
  input [18:0] Wgt_3_605, // sfix19_En18 
  input [18:0] Wgt_3_606, // sfix19_En18 
  input [18:0] Wgt_3_607, // sfix19_En18 
  input [18:0] Wgt_3_608, // sfix19_En18 
  input [18:0] Wgt_3_609, // sfix19_En18 
  input [18:0] Wgt_3_610, // sfix19_En18 
  input [18:0] Wgt_3_611, // sfix19_En18 
  input [18:0] Wgt_3_612, // sfix19_En18 
  input [18:0] Wgt_3_613, // sfix19_En18 
  input [18:0] Wgt_3_614, // sfix19_En18 
  input [18:0] Wgt_3_615, // sfix19_En18 
  input [18:0] Wgt_3_616, // sfix19_En18 
  input [18:0] Wgt_3_617, // sfix19_En18 
  input [18:0] Wgt_3_618, // sfix19_En18 
  input [18:0] Wgt_3_619, // sfix19_En18 
  input [18:0] Wgt_3_620, // sfix19_En18 
  input [18:0] Wgt_3_621, // sfix19_En18 
  input [18:0] Wgt_3_622, // sfix19_En18 
  input [18:0] Wgt_3_623, // sfix19_En18 
  input [18:0] Wgt_3_624, // sfix19_En18 
  input [18:0] Wgt_3_625, // sfix19_En18 
  input [18:0] Wgt_3_626, // sfix19_En18 
  input [18:0] Wgt_3_627, // sfix19_En18 
  input [18:0] Wgt_3_628, // sfix19_En18 
  input [18:0] Wgt_3_629, // sfix19_En18 
  input [18:0] Wgt_3_630, // sfix19_En18 
  input [18:0] Wgt_3_631, // sfix19_En18 
  input [18:0] Wgt_3_632, // sfix19_En18 
  input [18:0] Wgt_3_633, // sfix19_En18 
  input [18:0] Wgt_3_634, // sfix19_En18 
  input [18:0] Wgt_3_635, // sfix19_En18 
  input [18:0] Wgt_3_636, // sfix19_En18 
  input [18:0] Wgt_3_637, // sfix19_En18 
  input [18:0] Wgt_3_638, // sfix19_En18 
  input [18:0] Wgt_3_639, // sfix19_En18 
  input [18:0] Wgt_3_640, // sfix19_En18 
  input [18:0] Wgt_3_641, // sfix19_En18 
  input [18:0] Wgt_3_642, // sfix19_En18 
  input [18:0] Wgt_3_643, // sfix19_En18 
  input [18:0] Wgt_3_644, // sfix19_En18 
  input [18:0] Wgt_3_645, // sfix19_En18 
  input [18:0] Wgt_3_646, // sfix19_En18 
  input [18:0] Wgt_3_647, // sfix19_En18 
  input [18:0] Wgt_3_648, // sfix19_En18 
  input [18:0] Wgt_3_649, // sfix19_En18 
  input [18:0] Wgt_3_650, // sfix19_En18 
  input [18:0] Wgt_3_651, // sfix19_En18 
  input [18:0] Wgt_3_652, // sfix19_En18 
  input [18:0] Wgt_3_653, // sfix19_En18 
  input [18:0] Wgt_3_654, // sfix19_En18 
  input [18:0] Wgt_3_655, // sfix19_En18 
  input [18:0] Wgt_3_656, // sfix19_En18 
  input [18:0] Wgt_3_657, // sfix19_En18 
  input [18:0] Wgt_3_658, // sfix19_En18 
  input [18:0] Wgt_3_659, // sfix19_En18 
  input [18:0] Wgt_3_660, // sfix19_En18 
  input [18:0] Wgt_3_661, // sfix19_En18 
  input [18:0] Wgt_3_662, // sfix19_En18 
  input [18:0] Wgt_3_663, // sfix19_En18 
  input [18:0] Wgt_3_664, // sfix19_En18 
  input [18:0] Wgt_3_665, // sfix19_En18 
  input [18:0] Wgt_3_666, // sfix19_En18 
  input [18:0] Wgt_3_667, // sfix19_En18 
  input [18:0] Wgt_3_668, // sfix19_En18 
  input [18:0] Wgt_3_669, // sfix19_En18 
  input [18:0] Wgt_3_670, // sfix19_En18 
  input [18:0] Wgt_3_671, // sfix19_En18 
  input [18:0] Wgt_3_672, // sfix19_En18 
  input [18:0] Wgt_3_673, // sfix19_En18 
  input [18:0] Wgt_3_674, // sfix19_En18 
  input [18:0] Wgt_3_675, // sfix19_En18 
  input [18:0] Wgt_3_676, // sfix19_En18 
  input [18:0] Wgt_3_677, // sfix19_En18 
  input [18:0] Wgt_3_678, // sfix19_En18 
  input [18:0] Wgt_3_679, // sfix19_En18 
  input [18:0] Wgt_3_680, // sfix19_En18 
  input [18:0] Wgt_3_681, // sfix19_En18 
  input [18:0] Wgt_3_682, // sfix19_En18 
  input [18:0] Wgt_3_683, // sfix19_En18 
  input [18:0] Wgt_3_684, // sfix19_En18 
  input [18:0] Wgt_3_685, // sfix19_En18 
  input [18:0] Wgt_3_686, // sfix19_En18 
  input [18:0] Wgt_3_687, // sfix19_En18 
  input [18:0] Wgt_3_688, // sfix19_En18 
  input [18:0] Wgt_3_689, // sfix19_En18 
  input [18:0] Wgt_3_690, // sfix19_En18 
  input [18:0] Wgt_3_691, // sfix19_En18 
  input [18:0] Wgt_3_692, // sfix19_En18 
  input [18:0] Wgt_3_693, // sfix19_En18 
  input [18:0] Wgt_3_694, // sfix19_En18 
  input [18:0] Wgt_3_695, // sfix19_En18 
  input [18:0] Wgt_3_696, // sfix19_En18 
  input [18:0] Wgt_3_697, // sfix19_En18 
  input [18:0] Wgt_3_698, // sfix19_En18 
  input [18:0] Wgt_3_699, // sfix19_En18 
  input [18:0] Wgt_3_700, // sfix19_En18 
  input [18:0] Wgt_3_701, // sfix19_En18 
  input [18:0] Wgt_3_702, // sfix19_En18 
  input [18:0] Wgt_3_703, // sfix19_En18 
  input [18:0] Wgt_3_704, // sfix19_En18 
  input [18:0] Wgt_3_705, // sfix19_En18 
  input [18:0] Wgt_3_706, // sfix19_En18 
  input [18:0] Wgt_3_707, // sfix19_En18 
  input [18:0] Wgt_3_708, // sfix19_En18 
  input [18:0] Wgt_3_709, // sfix19_En18 
  input [18:0] Wgt_3_710, // sfix19_En18 
  input [18:0] Wgt_3_711, // sfix19_En18 
  input [18:0] Wgt_3_712, // sfix19_En18 
  input [18:0] Wgt_3_713, // sfix19_En18 
  input [18:0] Wgt_3_714, // sfix19_En18 
  input [18:0] Wgt_3_715, // sfix19_En18 
  input [18:0] Wgt_3_716, // sfix19_En18 
  input [18:0] Wgt_3_717, // sfix19_En18 
  input [18:0] Wgt_3_718, // sfix19_En18 
  input [18:0] Wgt_3_719, // sfix19_En18 
  input [18:0] Wgt_3_720, // sfix19_En18 
  input [18:0] Wgt_3_721, // sfix19_En18 
  input [18:0] Wgt_3_722, // sfix19_En18 
  input [18:0] Wgt_3_723, // sfix19_En18 
  input [18:0] Wgt_3_724, // sfix19_En18 
  input [18:0] Wgt_3_725, // sfix19_En18 
  input [18:0] Wgt_3_726, // sfix19_En18 
  input [18:0] Wgt_3_727, // sfix19_En18 
  input [18:0] Wgt_3_728, // sfix19_En18 
  input [18:0] Wgt_3_729, // sfix19_En18 
  input [18:0] Wgt_3_730, // sfix19_En18 
  input [18:0] Wgt_3_731, // sfix19_En18 
  input [18:0] Wgt_3_732, // sfix19_En18 
  input [18:0] Wgt_3_733, // sfix19_En18 
  input [18:0] Wgt_3_734, // sfix19_En18 
  input [18:0] Wgt_3_735, // sfix19_En18 
  input [18:0] Wgt_3_736, // sfix19_En18 
  input [18:0] Wgt_3_737, // sfix19_En18 
  input [18:0] Wgt_3_738, // sfix19_En18 
  input [18:0] Wgt_3_739, // sfix19_En18 
  input [18:0] Wgt_3_740, // sfix19_En18 
  input [18:0] Wgt_3_741, // sfix19_En18 
  input [18:0] Wgt_3_742, // sfix19_En18 
  input [18:0] Wgt_3_743, // sfix19_En18 
  input [18:0] Wgt_3_744, // sfix19_En18 
  input [18:0] Wgt_3_745, // sfix19_En18 
  input [18:0] Wgt_3_746, // sfix19_En18 
  input [18:0] Wgt_3_747, // sfix19_En18 
  input [18:0] Wgt_3_748, // sfix19_En18 
  input [18:0] Wgt_3_749, // sfix19_En18 
  input [18:0] Wgt_3_750, // sfix19_En18 
  input [18:0] Wgt_3_751, // sfix19_En18 
  input [18:0] Wgt_3_752, // sfix19_En18 
  input [18:0] Wgt_3_753, // sfix19_En18 
  input [18:0] Wgt_3_754, // sfix19_En18 
  input [18:0] Wgt_3_755, // sfix19_En18 
  input [18:0] Wgt_3_756, // sfix19_En18 
  input [18:0] Wgt_3_757, // sfix19_En18 
  input [18:0] Wgt_3_758, // sfix19_En18 
  input [18:0] Wgt_3_759, // sfix19_En18 
  input [18:0] Wgt_3_760, // sfix19_En18 
  input [18:0] Wgt_3_761, // sfix19_En18 
  input [18:0] Wgt_3_762, // sfix19_En18 
  input [18:0] Wgt_3_763, // sfix19_En18 
  input [18:0] Wgt_3_764, // sfix19_En18 
  input [18:0] Wgt_3_765, // sfix19_En18 
  input [18:0] Wgt_3_766, // sfix19_En18 
  input [18:0] Wgt_3_767, // sfix19_En18 
  input [18:0] Wgt_3_768, // sfix19_En18 
  input [18:0] Wgt_3_769, // sfix19_En18 
  input [18:0] Wgt_3_770, // sfix19_En18 
  input [18:0] Wgt_3_771, // sfix19_En18 
  input [18:0] Wgt_3_772, // sfix19_En18 
  input [18:0] Wgt_3_773, // sfix19_En18 
  input [18:0] Wgt_3_774, // sfix19_En18 
  input [18:0] Wgt_3_775, // sfix19_En18 
  input [18:0] Wgt_3_776, // sfix19_En18 
  input [18:0] Wgt_3_777, // sfix19_En18 
  input [18:0] Wgt_3_778, // sfix19_En18 
  input [18:0] Wgt_3_779, // sfix19_En18 
  input [18:0] Wgt_3_780, // sfix19_En18 
  input [18:0] Wgt_3_781, // sfix19_En18 
  input [18:0] Wgt_3_782, // sfix19_En18 
  input [18:0] Wgt_3_783, // sfix19_En18 
  input [18:0] Wgt_3_784, // sfix19_En18 
  input [18:0] Wgt_4_0, // sfix19_En18 
  input [18:0] Wgt_4_1, // sfix19_En18 
  input [18:0] Wgt_4_2, // sfix19_En18 
  input [18:0] Wgt_4_3, // sfix19_En18 
  input [18:0] Wgt_4_4, // sfix19_En18 
  input [18:0] Wgt_4_5, // sfix19_En18 
  input [18:0] Wgt_4_6, // sfix19_En18 
  input [18:0] Wgt_4_7, // sfix19_En18 
  input [18:0] Wgt_4_8, // sfix19_En18 
  input [18:0] Wgt_4_9, // sfix19_En18 
  input [18:0] Wgt_4_10, // sfix19_En18 
  input [18:0] Wgt_4_11, // sfix19_En18 
  input [18:0] Wgt_4_12, // sfix19_En18 
  input [18:0] Wgt_4_13, // sfix19_En18 
  input [18:0] Wgt_4_14, // sfix19_En18 
  input [18:0] Wgt_4_15, // sfix19_En18 
  input [18:0] Wgt_4_16, // sfix19_En18 
  input [18:0] Wgt_4_17, // sfix19_En18 
  input [18:0] Wgt_4_18, // sfix19_En18 
  input [18:0] Wgt_4_19, // sfix19_En18 
  input [18:0] Wgt_4_20, // sfix19_En18 
  input [18:0] Wgt_4_21, // sfix19_En18 
  input [18:0] Wgt_4_22, // sfix19_En18 
  input [18:0] Wgt_4_23, // sfix19_En18 
  input [18:0] Wgt_4_24, // sfix19_En18 
  input [18:0] Wgt_4_25, // sfix19_En18 
  input [18:0] Wgt_4_26, // sfix19_En18 
  input [18:0] Wgt_4_27, // sfix19_En18 
  input [18:0] Wgt_4_28, // sfix19_En18 
  input [18:0] Wgt_4_29, // sfix19_En18 
  input [18:0] Wgt_4_30, // sfix19_En18 
  input [18:0] Wgt_4_31, // sfix19_En18 
  input [18:0] Wgt_4_32, // sfix19_En18 
  input [18:0] Wgt_4_33, // sfix19_En18 
  input [18:0] Wgt_4_34, // sfix19_En18 
  input [18:0] Wgt_4_35, // sfix19_En18 
  input [18:0] Wgt_4_36, // sfix19_En18 
  input [18:0] Wgt_4_37, // sfix19_En18 
  input [18:0] Wgt_4_38, // sfix19_En18 
  input [18:0] Wgt_4_39, // sfix19_En18 
  input [18:0] Wgt_4_40, // sfix19_En18 
  input [18:0] Wgt_4_41, // sfix19_En18 
  input [18:0] Wgt_4_42, // sfix19_En18 
  input [18:0] Wgt_4_43, // sfix19_En18 
  input [18:0] Wgt_4_44, // sfix19_En18 
  input [18:0] Wgt_4_45, // sfix19_En18 
  input [18:0] Wgt_4_46, // sfix19_En18 
  input [18:0] Wgt_4_47, // sfix19_En18 
  input [18:0] Wgt_4_48, // sfix19_En18 
  input [18:0] Wgt_4_49, // sfix19_En18 
  input [18:0] Wgt_4_50, // sfix19_En18 
  input [18:0] Wgt_4_51, // sfix19_En18 
  input [18:0] Wgt_4_52, // sfix19_En18 
  input [18:0] Wgt_4_53, // sfix19_En18 
  input [18:0] Wgt_4_54, // sfix19_En18 
  input [18:0] Wgt_4_55, // sfix19_En18 
  input [18:0] Wgt_4_56, // sfix19_En18 
  input [18:0] Wgt_4_57, // sfix19_En18 
  input [18:0] Wgt_4_58, // sfix19_En18 
  input [18:0] Wgt_4_59, // sfix19_En18 
  input [18:0] Wgt_4_60, // sfix19_En18 
  input [18:0] Wgt_4_61, // sfix19_En18 
  input [18:0] Wgt_4_62, // sfix19_En18 
  input [18:0] Wgt_4_63, // sfix19_En18 
  input [18:0] Wgt_4_64, // sfix19_En18 
  input [18:0] Wgt_4_65, // sfix19_En18 
  input [18:0] Wgt_4_66, // sfix19_En18 
  input [18:0] Wgt_4_67, // sfix19_En18 
  input [18:0] Wgt_4_68, // sfix19_En18 
  input [18:0] Wgt_4_69, // sfix19_En18 
  input [18:0] Wgt_4_70, // sfix19_En18 
  input [18:0] Wgt_4_71, // sfix19_En18 
  input [18:0] Wgt_4_72, // sfix19_En18 
  input [18:0] Wgt_4_73, // sfix19_En18 
  input [18:0] Wgt_4_74, // sfix19_En18 
  input [18:0] Wgt_4_75, // sfix19_En18 
  input [18:0] Wgt_4_76, // sfix19_En18 
  input [18:0] Wgt_4_77, // sfix19_En18 
  input [18:0] Wgt_4_78, // sfix19_En18 
  input [18:0] Wgt_4_79, // sfix19_En18 
  input [18:0] Wgt_4_80, // sfix19_En18 
  input [18:0] Wgt_4_81, // sfix19_En18 
  input [18:0] Wgt_4_82, // sfix19_En18 
  input [18:0] Wgt_4_83, // sfix19_En18 
  input [18:0] Wgt_4_84, // sfix19_En18 
  input [18:0] Wgt_4_85, // sfix19_En18 
  input [18:0] Wgt_4_86, // sfix19_En18 
  input [18:0] Wgt_4_87, // sfix19_En18 
  input [18:0] Wgt_4_88, // sfix19_En18 
  input [18:0] Wgt_4_89, // sfix19_En18 
  input [18:0] Wgt_4_90, // sfix19_En18 
  input [18:0] Wgt_4_91, // sfix19_En18 
  input [18:0] Wgt_4_92, // sfix19_En18 
  input [18:0] Wgt_4_93, // sfix19_En18 
  input [18:0] Wgt_4_94, // sfix19_En18 
  input [18:0] Wgt_4_95, // sfix19_En18 
  input [18:0] Wgt_4_96, // sfix19_En18 
  input [18:0] Wgt_4_97, // sfix19_En18 
  input [18:0] Wgt_4_98, // sfix19_En18 
  input [18:0] Wgt_4_99, // sfix19_En18 
  input [18:0] Wgt_4_100, // sfix19_En18 
  input [18:0] Wgt_4_101, // sfix19_En18 
  input [18:0] Wgt_4_102, // sfix19_En18 
  input [18:0] Wgt_4_103, // sfix19_En18 
  input [18:0] Wgt_4_104, // sfix19_En18 
  input [18:0] Wgt_4_105, // sfix19_En18 
  input [18:0] Wgt_4_106, // sfix19_En18 
  input [18:0] Wgt_4_107, // sfix19_En18 
  input [18:0] Wgt_4_108, // sfix19_En18 
  input [18:0] Wgt_4_109, // sfix19_En18 
  input [18:0] Wgt_4_110, // sfix19_En18 
  input [18:0] Wgt_4_111, // sfix19_En18 
  input [18:0] Wgt_4_112, // sfix19_En18 
  input [18:0] Wgt_4_113, // sfix19_En18 
  input [18:0] Wgt_4_114, // sfix19_En18 
  input [18:0] Wgt_4_115, // sfix19_En18 
  input [18:0] Wgt_4_116, // sfix19_En18 
  input [18:0] Wgt_4_117, // sfix19_En18 
  input [18:0] Wgt_4_118, // sfix19_En18 
  input [18:0] Wgt_4_119, // sfix19_En18 
  input [18:0] Wgt_4_120, // sfix19_En18 
  input [18:0] Wgt_4_121, // sfix19_En18 
  input [18:0] Wgt_4_122, // sfix19_En18 
  input [18:0] Wgt_4_123, // sfix19_En18 
  input [18:0] Wgt_4_124, // sfix19_En18 
  input [18:0] Wgt_4_125, // sfix19_En18 
  input [18:0] Wgt_4_126, // sfix19_En18 
  input [18:0] Wgt_4_127, // sfix19_En18 
  input [18:0] Wgt_4_128, // sfix19_En18 
  input [18:0] Wgt_4_129, // sfix19_En18 
  input [18:0] Wgt_4_130, // sfix19_En18 
  input [18:0] Wgt_4_131, // sfix19_En18 
  input [18:0] Wgt_4_132, // sfix19_En18 
  input [18:0] Wgt_4_133, // sfix19_En18 
  input [18:0] Wgt_4_134, // sfix19_En18 
  input [18:0] Wgt_4_135, // sfix19_En18 
  input [18:0] Wgt_4_136, // sfix19_En18 
  input [18:0] Wgt_4_137, // sfix19_En18 
  input [18:0] Wgt_4_138, // sfix19_En18 
  input [18:0] Wgt_4_139, // sfix19_En18 
  input [18:0] Wgt_4_140, // sfix19_En18 
  input [18:0] Wgt_4_141, // sfix19_En18 
  input [18:0] Wgt_4_142, // sfix19_En18 
  input [18:0] Wgt_4_143, // sfix19_En18 
  input [18:0] Wgt_4_144, // sfix19_En18 
  input [18:0] Wgt_4_145, // sfix19_En18 
  input [18:0] Wgt_4_146, // sfix19_En18 
  input [18:0] Wgt_4_147, // sfix19_En18 
  input [18:0] Wgt_4_148, // sfix19_En18 
  input [18:0] Wgt_4_149, // sfix19_En18 
  input [18:0] Wgt_4_150, // sfix19_En18 
  input [18:0] Wgt_4_151, // sfix19_En18 
  input [18:0] Wgt_4_152, // sfix19_En18 
  input [18:0] Wgt_4_153, // sfix19_En18 
  input [18:0] Wgt_4_154, // sfix19_En18 
  input [18:0] Wgt_4_155, // sfix19_En18 
  input [18:0] Wgt_4_156, // sfix19_En18 
  input [18:0] Wgt_4_157, // sfix19_En18 
  input [18:0] Wgt_4_158, // sfix19_En18 
  input [18:0] Wgt_4_159, // sfix19_En18 
  input [18:0] Wgt_4_160, // sfix19_En18 
  input [18:0] Wgt_4_161, // sfix19_En18 
  input [18:0] Wgt_4_162, // sfix19_En18 
  input [18:0] Wgt_4_163, // sfix19_En18 
  input [18:0] Wgt_4_164, // sfix19_En18 
  input [18:0] Wgt_4_165, // sfix19_En18 
  input [18:0] Wgt_4_166, // sfix19_En18 
  input [18:0] Wgt_4_167, // sfix19_En18 
  input [18:0] Wgt_4_168, // sfix19_En18 
  input [18:0] Wgt_4_169, // sfix19_En18 
  input [18:0] Wgt_4_170, // sfix19_En18 
  input [18:0] Wgt_4_171, // sfix19_En18 
  input [18:0] Wgt_4_172, // sfix19_En18 
  input [18:0] Wgt_4_173, // sfix19_En18 
  input [18:0] Wgt_4_174, // sfix19_En18 
  input [18:0] Wgt_4_175, // sfix19_En18 
  input [18:0] Wgt_4_176, // sfix19_En18 
  input [18:0] Wgt_4_177, // sfix19_En18 
  input [18:0] Wgt_4_178, // sfix19_En18 
  input [18:0] Wgt_4_179, // sfix19_En18 
  input [18:0] Wgt_4_180, // sfix19_En18 
  input [18:0] Wgt_4_181, // sfix19_En18 
  input [18:0] Wgt_4_182, // sfix19_En18 
  input [18:0] Wgt_4_183, // sfix19_En18 
  input [18:0] Wgt_4_184, // sfix19_En18 
  input [18:0] Wgt_4_185, // sfix19_En18 
  input [18:0] Wgt_4_186, // sfix19_En18 
  input [18:0] Wgt_4_187, // sfix19_En18 
  input [18:0] Wgt_4_188, // sfix19_En18 
  input [18:0] Wgt_4_189, // sfix19_En18 
  input [18:0] Wgt_4_190, // sfix19_En18 
  input [18:0] Wgt_4_191, // sfix19_En18 
  input [18:0] Wgt_4_192, // sfix19_En18 
  input [18:0] Wgt_4_193, // sfix19_En18 
  input [18:0] Wgt_4_194, // sfix19_En18 
  input [18:0] Wgt_4_195, // sfix19_En18 
  input [18:0] Wgt_4_196, // sfix19_En18 
  input [18:0] Wgt_4_197, // sfix19_En18 
  input [18:0] Wgt_4_198, // sfix19_En18 
  input [18:0] Wgt_4_199, // sfix19_En18 
  input [18:0] Wgt_4_200, // sfix19_En18 
  input [18:0] Wgt_4_201, // sfix19_En18 
  input [18:0] Wgt_4_202, // sfix19_En18 
  input [18:0] Wgt_4_203, // sfix19_En18 
  input [18:0] Wgt_4_204, // sfix19_En18 
  input [18:0] Wgt_4_205, // sfix19_En18 
  input [18:0] Wgt_4_206, // sfix19_En18 
  input [18:0] Wgt_4_207, // sfix19_En18 
  input [18:0] Wgt_4_208, // sfix19_En18 
  input [18:0] Wgt_4_209, // sfix19_En18 
  input [18:0] Wgt_4_210, // sfix19_En18 
  input [18:0] Wgt_4_211, // sfix19_En18 
  input [18:0] Wgt_4_212, // sfix19_En18 
  input [18:0] Wgt_4_213, // sfix19_En18 
  input [18:0] Wgt_4_214, // sfix19_En18 
  input [18:0] Wgt_4_215, // sfix19_En18 
  input [18:0] Wgt_4_216, // sfix19_En18 
  input [18:0] Wgt_4_217, // sfix19_En18 
  input [18:0] Wgt_4_218, // sfix19_En18 
  input [18:0] Wgt_4_219, // sfix19_En18 
  input [18:0] Wgt_4_220, // sfix19_En18 
  input [18:0] Wgt_4_221, // sfix19_En18 
  input [18:0] Wgt_4_222, // sfix19_En18 
  input [18:0] Wgt_4_223, // sfix19_En18 
  input [18:0] Wgt_4_224, // sfix19_En18 
  input [18:0] Wgt_4_225, // sfix19_En18 
  input [18:0] Wgt_4_226, // sfix19_En18 
  input [18:0] Wgt_4_227, // sfix19_En18 
  input [18:0] Wgt_4_228, // sfix19_En18 
  input [18:0] Wgt_4_229, // sfix19_En18 
  input [18:0] Wgt_4_230, // sfix19_En18 
  input [18:0] Wgt_4_231, // sfix19_En18 
  input [18:0] Wgt_4_232, // sfix19_En18 
  input [18:0] Wgt_4_233, // sfix19_En18 
  input [18:0] Wgt_4_234, // sfix19_En18 
  input [18:0] Wgt_4_235, // sfix19_En18 
  input [18:0] Wgt_4_236, // sfix19_En18 
  input [18:0] Wgt_4_237, // sfix19_En18 
  input [18:0] Wgt_4_238, // sfix19_En18 
  input [18:0] Wgt_4_239, // sfix19_En18 
  input [18:0] Wgt_4_240, // sfix19_En18 
  input [18:0] Wgt_4_241, // sfix19_En18 
  input [18:0] Wgt_4_242, // sfix19_En18 
  input [18:0] Wgt_4_243, // sfix19_En18 
  input [18:0] Wgt_4_244, // sfix19_En18 
  input [18:0] Wgt_4_245, // sfix19_En18 
  input [18:0] Wgt_4_246, // sfix19_En18 
  input [18:0] Wgt_4_247, // sfix19_En18 
  input [18:0] Wgt_4_248, // sfix19_En18 
  input [18:0] Wgt_4_249, // sfix19_En18 
  input [18:0] Wgt_4_250, // sfix19_En18 
  input [18:0] Wgt_4_251, // sfix19_En18 
  input [18:0] Wgt_4_252, // sfix19_En18 
  input [18:0] Wgt_4_253, // sfix19_En18 
  input [18:0] Wgt_4_254, // sfix19_En18 
  input [18:0] Wgt_4_255, // sfix19_En18 
  input [18:0] Wgt_4_256, // sfix19_En18 
  input [18:0] Wgt_4_257, // sfix19_En18 
  input [18:0] Wgt_4_258, // sfix19_En18 
  input [18:0] Wgt_4_259, // sfix19_En18 
  input [18:0] Wgt_4_260, // sfix19_En18 
  input [18:0] Wgt_4_261, // sfix19_En18 
  input [18:0] Wgt_4_262, // sfix19_En18 
  input [18:0] Wgt_4_263, // sfix19_En18 
  input [18:0] Wgt_4_264, // sfix19_En18 
  input [18:0] Wgt_4_265, // sfix19_En18 
  input [18:0] Wgt_4_266, // sfix19_En18 
  input [18:0] Wgt_4_267, // sfix19_En18 
  input [18:0] Wgt_4_268, // sfix19_En18 
  input [18:0] Wgt_4_269, // sfix19_En18 
  input [18:0] Wgt_4_270, // sfix19_En18 
  input [18:0] Wgt_4_271, // sfix19_En18 
  input [18:0] Wgt_4_272, // sfix19_En18 
  input [18:0] Wgt_4_273, // sfix19_En18 
  input [18:0] Wgt_4_274, // sfix19_En18 
  input [18:0] Wgt_4_275, // sfix19_En18 
  input [18:0] Wgt_4_276, // sfix19_En18 
  input [18:0] Wgt_4_277, // sfix19_En18 
  input [18:0] Wgt_4_278, // sfix19_En18 
  input [18:0] Wgt_4_279, // sfix19_En18 
  input [18:0] Wgt_4_280, // sfix19_En18 
  input [18:0] Wgt_4_281, // sfix19_En18 
  input [18:0] Wgt_4_282, // sfix19_En18 
  input [18:0] Wgt_4_283, // sfix19_En18 
  input [18:0] Wgt_4_284, // sfix19_En18 
  input [18:0] Wgt_4_285, // sfix19_En18 
  input [18:0] Wgt_4_286, // sfix19_En18 
  input [18:0] Wgt_4_287, // sfix19_En18 
  input [18:0] Wgt_4_288, // sfix19_En18 
  input [18:0] Wgt_4_289, // sfix19_En18 
  input [18:0] Wgt_4_290, // sfix19_En18 
  input [18:0] Wgt_4_291, // sfix19_En18 
  input [18:0] Wgt_4_292, // sfix19_En18 
  input [18:0] Wgt_4_293, // sfix19_En18 
  input [18:0] Wgt_4_294, // sfix19_En18 
  input [18:0] Wgt_4_295, // sfix19_En18 
  input [18:0] Wgt_4_296, // sfix19_En18 
  input [18:0] Wgt_4_297, // sfix19_En18 
  input [18:0] Wgt_4_298, // sfix19_En18 
  input [18:0] Wgt_4_299, // sfix19_En18 
  input [18:0] Wgt_4_300, // sfix19_En18 
  input [18:0] Wgt_4_301, // sfix19_En18 
  input [18:0] Wgt_4_302, // sfix19_En18 
  input [18:0] Wgt_4_303, // sfix19_En18 
  input [18:0] Wgt_4_304, // sfix19_En18 
  input [18:0] Wgt_4_305, // sfix19_En18 
  input [18:0] Wgt_4_306, // sfix19_En18 
  input [18:0] Wgt_4_307, // sfix19_En18 
  input [18:0] Wgt_4_308, // sfix19_En18 
  input [18:0] Wgt_4_309, // sfix19_En18 
  input [18:0] Wgt_4_310, // sfix19_En18 
  input [18:0] Wgt_4_311, // sfix19_En18 
  input [18:0] Wgt_4_312, // sfix19_En18 
  input [18:0] Wgt_4_313, // sfix19_En18 
  input [18:0] Wgt_4_314, // sfix19_En18 
  input [18:0] Wgt_4_315, // sfix19_En18 
  input [18:0] Wgt_4_316, // sfix19_En18 
  input [18:0] Wgt_4_317, // sfix19_En18 
  input [18:0] Wgt_4_318, // sfix19_En18 
  input [18:0] Wgt_4_319, // sfix19_En18 
  input [18:0] Wgt_4_320, // sfix19_En18 
  input [18:0] Wgt_4_321, // sfix19_En18 
  input [18:0] Wgt_4_322, // sfix19_En18 
  input [18:0] Wgt_4_323, // sfix19_En18 
  input [18:0] Wgt_4_324, // sfix19_En18 
  input [18:0] Wgt_4_325, // sfix19_En18 
  input [18:0] Wgt_4_326, // sfix19_En18 
  input [18:0] Wgt_4_327, // sfix19_En18 
  input [18:0] Wgt_4_328, // sfix19_En18 
  input [18:0] Wgt_4_329, // sfix19_En18 
  input [18:0] Wgt_4_330, // sfix19_En18 
  input [18:0] Wgt_4_331, // sfix19_En18 
  input [18:0] Wgt_4_332, // sfix19_En18 
  input [18:0] Wgt_4_333, // sfix19_En18 
  input [18:0] Wgt_4_334, // sfix19_En18 
  input [18:0] Wgt_4_335, // sfix19_En18 
  input [18:0] Wgt_4_336, // sfix19_En18 
  input [18:0] Wgt_4_337, // sfix19_En18 
  input [18:0] Wgt_4_338, // sfix19_En18 
  input [18:0] Wgt_4_339, // sfix19_En18 
  input [18:0] Wgt_4_340, // sfix19_En18 
  input [18:0] Wgt_4_341, // sfix19_En18 
  input [18:0] Wgt_4_342, // sfix19_En18 
  input [18:0] Wgt_4_343, // sfix19_En18 
  input [18:0] Wgt_4_344, // sfix19_En18 
  input [18:0] Wgt_4_345, // sfix19_En18 
  input [18:0] Wgt_4_346, // sfix19_En18 
  input [18:0] Wgt_4_347, // sfix19_En18 
  input [18:0] Wgt_4_348, // sfix19_En18 
  input [18:0] Wgt_4_349, // sfix19_En18 
  input [18:0] Wgt_4_350, // sfix19_En18 
  input [18:0] Wgt_4_351, // sfix19_En18 
  input [18:0] Wgt_4_352, // sfix19_En18 
  input [18:0] Wgt_4_353, // sfix19_En18 
  input [18:0] Wgt_4_354, // sfix19_En18 
  input [18:0] Wgt_4_355, // sfix19_En18 
  input [18:0] Wgt_4_356, // sfix19_En18 
  input [18:0] Wgt_4_357, // sfix19_En18 
  input [18:0] Wgt_4_358, // sfix19_En18 
  input [18:0] Wgt_4_359, // sfix19_En18 
  input [18:0] Wgt_4_360, // sfix19_En18 
  input [18:0] Wgt_4_361, // sfix19_En18 
  input [18:0] Wgt_4_362, // sfix19_En18 
  input [18:0] Wgt_4_363, // sfix19_En18 
  input [18:0] Wgt_4_364, // sfix19_En18 
  input [18:0] Wgt_4_365, // sfix19_En18 
  input [18:0] Wgt_4_366, // sfix19_En18 
  input [18:0] Wgt_4_367, // sfix19_En18 
  input [18:0] Wgt_4_368, // sfix19_En18 
  input [18:0] Wgt_4_369, // sfix19_En18 
  input [18:0] Wgt_4_370, // sfix19_En18 
  input [18:0] Wgt_4_371, // sfix19_En18 
  input [18:0] Wgt_4_372, // sfix19_En18 
  input [18:0] Wgt_4_373, // sfix19_En18 
  input [18:0] Wgt_4_374, // sfix19_En18 
  input [18:0] Wgt_4_375, // sfix19_En18 
  input [18:0] Wgt_4_376, // sfix19_En18 
  input [18:0] Wgt_4_377, // sfix19_En18 
  input [18:0] Wgt_4_378, // sfix19_En18 
  input [18:0] Wgt_4_379, // sfix19_En18 
  input [18:0] Wgt_4_380, // sfix19_En18 
  input [18:0] Wgt_4_381, // sfix19_En18 
  input [18:0] Wgt_4_382, // sfix19_En18 
  input [18:0] Wgt_4_383, // sfix19_En18 
  input [18:0] Wgt_4_384, // sfix19_En18 
  input [18:0] Wgt_4_385, // sfix19_En18 
  input [18:0] Wgt_4_386, // sfix19_En18 
  input [18:0] Wgt_4_387, // sfix19_En18 
  input [18:0] Wgt_4_388, // sfix19_En18 
  input [18:0] Wgt_4_389, // sfix19_En18 
  input [18:0] Wgt_4_390, // sfix19_En18 
  input [18:0] Wgt_4_391, // sfix19_En18 
  input [18:0] Wgt_4_392, // sfix19_En18 
  input [18:0] Wgt_4_393, // sfix19_En18 
  input [18:0] Wgt_4_394, // sfix19_En18 
  input [18:0] Wgt_4_395, // sfix19_En18 
  input [18:0] Wgt_4_396, // sfix19_En18 
  input [18:0] Wgt_4_397, // sfix19_En18 
  input [18:0] Wgt_4_398, // sfix19_En18 
  input [18:0] Wgt_4_399, // sfix19_En18 
  input [18:0] Wgt_4_400, // sfix19_En18 
  input [18:0] Wgt_4_401, // sfix19_En18 
  input [18:0] Wgt_4_402, // sfix19_En18 
  input [18:0] Wgt_4_403, // sfix19_En18 
  input [18:0] Wgt_4_404, // sfix19_En18 
  input [18:0] Wgt_4_405, // sfix19_En18 
  input [18:0] Wgt_4_406, // sfix19_En18 
  input [18:0] Wgt_4_407, // sfix19_En18 
  input [18:0] Wgt_4_408, // sfix19_En18 
  input [18:0] Wgt_4_409, // sfix19_En18 
  input [18:0] Wgt_4_410, // sfix19_En18 
  input [18:0] Wgt_4_411, // sfix19_En18 
  input [18:0] Wgt_4_412, // sfix19_En18 
  input [18:0] Wgt_4_413, // sfix19_En18 
  input [18:0] Wgt_4_414, // sfix19_En18 
  input [18:0] Wgt_4_415, // sfix19_En18 
  input [18:0] Wgt_4_416, // sfix19_En18 
  input [18:0] Wgt_4_417, // sfix19_En18 
  input [18:0] Wgt_4_418, // sfix19_En18 
  input [18:0] Wgt_4_419, // sfix19_En18 
  input [18:0] Wgt_4_420, // sfix19_En18 
  input [18:0] Wgt_4_421, // sfix19_En18 
  input [18:0] Wgt_4_422, // sfix19_En18 
  input [18:0] Wgt_4_423, // sfix19_En18 
  input [18:0] Wgt_4_424, // sfix19_En18 
  input [18:0] Wgt_4_425, // sfix19_En18 
  input [18:0] Wgt_4_426, // sfix19_En18 
  input [18:0] Wgt_4_427, // sfix19_En18 
  input [18:0] Wgt_4_428, // sfix19_En18 
  input [18:0] Wgt_4_429, // sfix19_En18 
  input [18:0] Wgt_4_430, // sfix19_En18 
  input [18:0] Wgt_4_431, // sfix19_En18 
  input [18:0] Wgt_4_432, // sfix19_En18 
  input [18:0] Wgt_4_433, // sfix19_En18 
  input [18:0] Wgt_4_434, // sfix19_En18 
  input [18:0] Wgt_4_435, // sfix19_En18 
  input [18:0] Wgt_4_436, // sfix19_En18 
  input [18:0] Wgt_4_437, // sfix19_En18 
  input [18:0] Wgt_4_438, // sfix19_En18 
  input [18:0] Wgt_4_439, // sfix19_En18 
  input [18:0] Wgt_4_440, // sfix19_En18 
  input [18:0] Wgt_4_441, // sfix19_En18 
  input [18:0] Wgt_4_442, // sfix19_En18 
  input [18:0] Wgt_4_443, // sfix19_En18 
  input [18:0] Wgt_4_444, // sfix19_En18 
  input [18:0] Wgt_4_445, // sfix19_En18 
  input [18:0] Wgt_4_446, // sfix19_En18 
  input [18:0] Wgt_4_447, // sfix19_En18 
  input [18:0] Wgt_4_448, // sfix19_En18 
  input [18:0] Wgt_4_449, // sfix19_En18 
  input [18:0] Wgt_4_450, // sfix19_En18 
  input [18:0] Wgt_4_451, // sfix19_En18 
  input [18:0] Wgt_4_452, // sfix19_En18 
  input [18:0] Wgt_4_453, // sfix19_En18 
  input [18:0] Wgt_4_454, // sfix19_En18 
  input [18:0] Wgt_4_455, // sfix19_En18 
  input [18:0] Wgt_4_456, // sfix19_En18 
  input [18:0] Wgt_4_457, // sfix19_En18 
  input [18:0] Wgt_4_458, // sfix19_En18 
  input [18:0] Wgt_4_459, // sfix19_En18 
  input [18:0] Wgt_4_460, // sfix19_En18 
  input [18:0] Wgt_4_461, // sfix19_En18 
  input [18:0] Wgt_4_462, // sfix19_En18 
  input [18:0] Wgt_4_463, // sfix19_En18 
  input [18:0] Wgt_4_464, // sfix19_En18 
  input [18:0] Wgt_4_465, // sfix19_En18 
  input [18:0] Wgt_4_466, // sfix19_En18 
  input [18:0] Wgt_4_467, // sfix19_En18 
  input [18:0] Wgt_4_468, // sfix19_En18 
  input [18:0] Wgt_4_469, // sfix19_En18 
  input [18:0] Wgt_4_470, // sfix19_En18 
  input [18:0] Wgt_4_471, // sfix19_En18 
  input [18:0] Wgt_4_472, // sfix19_En18 
  input [18:0] Wgt_4_473, // sfix19_En18 
  input [18:0] Wgt_4_474, // sfix19_En18 
  input [18:0] Wgt_4_475, // sfix19_En18 
  input [18:0] Wgt_4_476, // sfix19_En18 
  input [18:0] Wgt_4_477, // sfix19_En18 
  input [18:0] Wgt_4_478, // sfix19_En18 
  input [18:0] Wgt_4_479, // sfix19_En18 
  input [18:0] Wgt_4_480, // sfix19_En18 
  input [18:0] Wgt_4_481, // sfix19_En18 
  input [18:0] Wgt_4_482, // sfix19_En18 
  input [18:0] Wgt_4_483, // sfix19_En18 
  input [18:0] Wgt_4_484, // sfix19_En18 
  input [18:0] Wgt_4_485, // sfix19_En18 
  input [18:0] Wgt_4_486, // sfix19_En18 
  input [18:0] Wgt_4_487, // sfix19_En18 
  input [18:0] Wgt_4_488, // sfix19_En18 
  input [18:0] Wgt_4_489, // sfix19_En18 
  input [18:0] Wgt_4_490, // sfix19_En18 
  input [18:0] Wgt_4_491, // sfix19_En18 
  input [18:0] Wgt_4_492, // sfix19_En18 
  input [18:0] Wgt_4_493, // sfix19_En18 
  input [18:0] Wgt_4_494, // sfix19_En18 
  input [18:0] Wgt_4_495, // sfix19_En18 
  input [18:0] Wgt_4_496, // sfix19_En18 
  input [18:0] Wgt_4_497, // sfix19_En18 
  input [18:0] Wgt_4_498, // sfix19_En18 
  input [18:0] Wgt_4_499, // sfix19_En18 
  input [18:0] Wgt_4_500, // sfix19_En18 
  input [18:0] Wgt_4_501, // sfix19_En18 
  input [18:0] Wgt_4_502, // sfix19_En18 
  input [18:0] Wgt_4_503, // sfix19_En18 
  input [18:0] Wgt_4_504, // sfix19_En18 
  input [18:0] Wgt_4_505, // sfix19_En18 
  input [18:0] Wgt_4_506, // sfix19_En18 
  input [18:0] Wgt_4_507, // sfix19_En18 
  input [18:0] Wgt_4_508, // sfix19_En18 
  input [18:0] Wgt_4_509, // sfix19_En18 
  input [18:0] Wgt_4_510, // sfix19_En18 
  input [18:0] Wgt_4_511, // sfix19_En18 
  input [18:0] Wgt_4_512, // sfix19_En18 
  input [18:0] Wgt_4_513, // sfix19_En18 
  input [18:0] Wgt_4_514, // sfix19_En18 
  input [18:0] Wgt_4_515, // sfix19_En18 
  input [18:0] Wgt_4_516, // sfix19_En18 
  input [18:0] Wgt_4_517, // sfix19_En18 
  input [18:0] Wgt_4_518, // sfix19_En18 
  input [18:0] Wgt_4_519, // sfix19_En18 
  input [18:0] Wgt_4_520, // sfix19_En18 
  input [18:0] Wgt_4_521, // sfix19_En18 
  input [18:0] Wgt_4_522, // sfix19_En18 
  input [18:0] Wgt_4_523, // sfix19_En18 
  input [18:0] Wgt_4_524, // sfix19_En18 
  input [18:0] Wgt_4_525, // sfix19_En18 
  input [18:0] Wgt_4_526, // sfix19_En18 
  input [18:0] Wgt_4_527, // sfix19_En18 
  input [18:0] Wgt_4_528, // sfix19_En18 
  input [18:0] Wgt_4_529, // sfix19_En18 
  input [18:0] Wgt_4_530, // sfix19_En18 
  input [18:0] Wgt_4_531, // sfix19_En18 
  input [18:0] Wgt_4_532, // sfix19_En18 
  input [18:0] Wgt_4_533, // sfix19_En18 
  input [18:0] Wgt_4_534, // sfix19_En18 
  input [18:0] Wgt_4_535, // sfix19_En18 
  input [18:0] Wgt_4_536, // sfix19_En18 
  input [18:0] Wgt_4_537, // sfix19_En18 
  input [18:0] Wgt_4_538, // sfix19_En18 
  input [18:0] Wgt_4_539, // sfix19_En18 
  input [18:0] Wgt_4_540, // sfix19_En18 
  input [18:0] Wgt_4_541, // sfix19_En18 
  input [18:0] Wgt_4_542, // sfix19_En18 
  input [18:0] Wgt_4_543, // sfix19_En18 
  input [18:0] Wgt_4_544, // sfix19_En18 
  input [18:0] Wgt_4_545, // sfix19_En18 
  input [18:0] Wgt_4_546, // sfix19_En18 
  input [18:0] Wgt_4_547, // sfix19_En18 
  input [18:0] Wgt_4_548, // sfix19_En18 
  input [18:0] Wgt_4_549, // sfix19_En18 
  input [18:0] Wgt_4_550, // sfix19_En18 
  input [18:0] Wgt_4_551, // sfix19_En18 
  input [18:0] Wgt_4_552, // sfix19_En18 
  input [18:0] Wgt_4_553, // sfix19_En18 
  input [18:0] Wgt_4_554, // sfix19_En18 
  input [18:0] Wgt_4_555, // sfix19_En18 
  input [18:0] Wgt_4_556, // sfix19_En18 
  input [18:0] Wgt_4_557, // sfix19_En18 
  input [18:0] Wgt_4_558, // sfix19_En18 
  input [18:0] Wgt_4_559, // sfix19_En18 
  input [18:0] Wgt_4_560, // sfix19_En18 
  input [18:0] Wgt_4_561, // sfix19_En18 
  input [18:0] Wgt_4_562, // sfix19_En18 
  input [18:0] Wgt_4_563, // sfix19_En18 
  input [18:0] Wgt_4_564, // sfix19_En18 
  input [18:0] Wgt_4_565, // sfix19_En18 
  input [18:0] Wgt_4_566, // sfix19_En18 
  input [18:0] Wgt_4_567, // sfix19_En18 
  input [18:0] Wgt_4_568, // sfix19_En18 
  input [18:0] Wgt_4_569, // sfix19_En18 
  input [18:0] Wgt_4_570, // sfix19_En18 
  input [18:0] Wgt_4_571, // sfix19_En18 
  input [18:0] Wgt_4_572, // sfix19_En18 
  input [18:0] Wgt_4_573, // sfix19_En18 
  input [18:0] Wgt_4_574, // sfix19_En18 
  input [18:0] Wgt_4_575, // sfix19_En18 
  input [18:0] Wgt_4_576, // sfix19_En18 
  input [18:0] Wgt_4_577, // sfix19_En18 
  input [18:0] Wgt_4_578, // sfix19_En18 
  input [18:0] Wgt_4_579, // sfix19_En18 
  input [18:0] Wgt_4_580, // sfix19_En18 
  input [18:0] Wgt_4_581, // sfix19_En18 
  input [18:0] Wgt_4_582, // sfix19_En18 
  input [18:0] Wgt_4_583, // sfix19_En18 
  input [18:0] Wgt_4_584, // sfix19_En18 
  input [18:0] Wgt_4_585, // sfix19_En18 
  input [18:0] Wgt_4_586, // sfix19_En18 
  input [18:0] Wgt_4_587, // sfix19_En18 
  input [18:0] Wgt_4_588, // sfix19_En18 
  input [18:0] Wgt_4_589, // sfix19_En18 
  input [18:0] Wgt_4_590, // sfix19_En18 
  input [18:0] Wgt_4_591, // sfix19_En18 
  input [18:0] Wgt_4_592, // sfix19_En18 
  input [18:0] Wgt_4_593, // sfix19_En18 
  input [18:0] Wgt_4_594, // sfix19_En18 
  input [18:0] Wgt_4_595, // sfix19_En18 
  input [18:0] Wgt_4_596, // sfix19_En18 
  input [18:0] Wgt_4_597, // sfix19_En18 
  input [18:0] Wgt_4_598, // sfix19_En18 
  input [18:0] Wgt_4_599, // sfix19_En18 
  input [18:0] Wgt_4_600, // sfix19_En18 
  input [18:0] Wgt_4_601, // sfix19_En18 
  input [18:0] Wgt_4_602, // sfix19_En18 
  input [18:0] Wgt_4_603, // sfix19_En18 
  input [18:0] Wgt_4_604, // sfix19_En18 
  input [18:0] Wgt_4_605, // sfix19_En18 
  input [18:0] Wgt_4_606, // sfix19_En18 
  input [18:0] Wgt_4_607, // sfix19_En18 
  input [18:0] Wgt_4_608, // sfix19_En18 
  input [18:0] Wgt_4_609, // sfix19_En18 
  input [18:0] Wgt_4_610, // sfix19_En18 
  input [18:0] Wgt_4_611, // sfix19_En18 
  input [18:0] Wgt_4_612, // sfix19_En18 
  input [18:0] Wgt_4_613, // sfix19_En18 
  input [18:0] Wgt_4_614, // sfix19_En18 
  input [18:0] Wgt_4_615, // sfix19_En18 
  input [18:0] Wgt_4_616, // sfix19_En18 
  input [18:0] Wgt_4_617, // sfix19_En18 
  input [18:0] Wgt_4_618, // sfix19_En18 
  input [18:0] Wgt_4_619, // sfix19_En18 
  input [18:0] Wgt_4_620, // sfix19_En18 
  input [18:0] Wgt_4_621, // sfix19_En18 
  input [18:0] Wgt_4_622, // sfix19_En18 
  input [18:0] Wgt_4_623, // sfix19_En18 
  input [18:0] Wgt_4_624, // sfix19_En18 
  input [18:0] Wgt_4_625, // sfix19_En18 
  input [18:0] Wgt_4_626, // sfix19_En18 
  input [18:0] Wgt_4_627, // sfix19_En18 
  input [18:0] Wgt_4_628, // sfix19_En18 
  input [18:0] Wgt_4_629, // sfix19_En18 
  input [18:0] Wgt_4_630, // sfix19_En18 
  input [18:0] Wgt_4_631, // sfix19_En18 
  input [18:0] Wgt_4_632, // sfix19_En18 
  input [18:0] Wgt_4_633, // sfix19_En18 
  input [18:0] Wgt_4_634, // sfix19_En18 
  input [18:0] Wgt_4_635, // sfix19_En18 
  input [18:0] Wgt_4_636, // sfix19_En18 
  input [18:0] Wgt_4_637, // sfix19_En18 
  input [18:0] Wgt_4_638, // sfix19_En18 
  input [18:0] Wgt_4_639, // sfix19_En18 
  input [18:0] Wgt_4_640, // sfix19_En18 
  input [18:0] Wgt_4_641, // sfix19_En18 
  input [18:0] Wgt_4_642, // sfix19_En18 
  input [18:0] Wgt_4_643, // sfix19_En18 
  input [18:0] Wgt_4_644, // sfix19_En18 
  input [18:0] Wgt_4_645, // sfix19_En18 
  input [18:0] Wgt_4_646, // sfix19_En18 
  input [18:0] Wgt_4_647, // sfix19_En18 
  input [18:0] Wgt_4_648, // sfix19_En18 
  input [18:0] Wgt_4_649, // sfix19_En18 
  input [18:0] Wgt_4_650, // sfix19_En18 
  input [18:0] Wgt_4_651, // sfix19_En18 
  input [18:0] Wgt_4_652, // sfix19_En18 
  input [18:0] Wgt_4_653, // sfix19_En18 
  input [18:0] Wgt_4_654, // sfix19_En18 
  input [18:0] Wgt_4_655, // sfix19_En18 
  input [18:0] Wgt_4_656, // sfix19_En18 
  input [18:0] Wgt_4_657, // sfix19_En18 
  input [18:0] Wgt_4_658, // sfix19_En18 
  input [18:0] Wgt_4_659, // sfix19_En18 
  input [18:0] Wgt_4_660, // sfix19_En18 
  input [18:0] Wgt_4_661, // sfix19_En18 
  input [18:0] Wgt_4_662, // sfix19_En18 
  input [18:0] Wgt_4_663, // sfix19_En18 
  input [18:0] Wgt_4_664, // sfix19_En18 
  input [18:0] Wgt_4_665, // sfix19_En18 
  input [18:0] Wgt_4_666, // sfix19_En18 
  input [18:0] Wgt_4_667, // sfix19_En18 
  input [18:0] Wgt_4_668, // sfix19_En18 
  input [18:0] Wgt_4_669, // sfix19_En18 
  input [18:0] Wgt_4_670, // sfix19_En18 
  input [18:0] Wgt_4_671, // sfix19_En18 
  input [18:0] Wgt_4_672, // sfix19_En18 
  input [18:0] Wgt_4_673, // sfix19_En18 
  input [18:0] Wgt_4_674, // sfix19_En18 
  input [18:0] Wgt_4_675, // sfix19_En18 
  input [18:0] Wgt_4_676, // sfix19_En18 
  input [18:0] Wgt_4_677, // sfix19_En18 
  input [18:0] Wgt_4_678, // sfix19_En18 
  input [18:0] Wgt_4_679, // sfix19_En18 
  input [18:0] Wgt_4_680, // sfix19_En18 
  input [18:0] Wgt_4_681, // sfix19_En18 
  input [18:0] Wgt_4_682, // sfix19_En18 
  input [18:0] Wgt_4_683, // sfix19_En18 
  input [18:0] Wgt_4_684, // sfix19_En18 
  input [18:0] Wgt_4_685, // sfix19_En18 
  input [18:0] Wgt_4_686, // sfix19_En18 
  input [18:0] Wgt_4_687, // sfix19_En18 
  input [18:0] Wgt_4_688, // sfix19_En18 
  input [18:0] Wgt_4_689, // sfix19_En18 
  input [18:0] Wgt_4_690, // sfix19_En18 
  input [18:0] Wgt_4_691, // sfix19_En18 
  input [18:0] Wgt_4_692, // sfix19_En18 
  input [18:0] Wgt_4_693, // sfix19_En18 
  input [18:0] Wgt_4_694, // sfix19_En18 
  input [18:0] Wgt_4_695, // sfix19_En18 
  input [18:0] Wgt_4_696, // sfix19_En18 
  input [18:0] Wgt_4_697, // sfix19_En18 
  input [18:0] Wgt_4_698, // sfix19_En18 
  input [18:0] Wgt_4_699, // sfix19_En18 
  input [18:0] Wgt_4_700, // sfix19_En18 
  input [18:0] Wgt_4_701, // sfix19_En18 
  input [18:0] Wgt_4_702, // sfix19_En18 
  input [18:0] Wgt_4_703, // sfix19_En18 
  input [18:0] Wgt_4_704, // sfix19_En18 
  input [18:0] Wgt_4_705, // sfix19_En18 
  input [18:0] Wgt_4_706, // sfix19_En18 
  input [18:0] Wgt_4_707, // sfix19_En18 
  input [18:0] Wgt_4_708, // sfix19_En18 
  input [18:0] Wgt_4_709, // sfix19_En18 
  input [18:0] Wgt_4_710, // sfix19_En18 
  input [18:0] Wgt_4_711, // sfix19_En18 
  input [18:0] Wgt_4_712, // sfix19_En18 
  input [18:0] Wgt_4_713, // sfix19_En18 
  input [18:0] Wgt_4_714, // sfix19_En18 
  input [18:0] Wgt_4_715, // sfix19_En18 
  input [18:0] Wgt_4_716, // sfix19_En18 
  input [18:0] Wgt_4_717, // sfix19_En18 
  input [18:0] Wgt_4_718, // sfix19_En18 
  input [18:0] Wgt_4_719, // sfix19_En18 
  input [18:0] Wgt_4_720, // sfix19_En18 
  input [18:0] Wgt_4_721, // sfix19_En18 
  input [18:0] Wgt_4_722, // sfix19_En18 
  input [18:0] Wgt_4_723, // sfix19_En18 
  input [18:0] Wgt_4_724, // sfix19_En18 
  input [18:0] Wgt_4_725, // sfix19_En18 
  input [18:0] Wgt_4_726, // sfix19_En18 
  input [18:0] Wgt_4_727, // sfix19_En18 
  input [18:0] Wgt_4_728, // sfix19_En18 
  input [18:0] Wgt_4_729, // sfix19_En18 
  input [18:0] Wgt_4_730, // sfix19_En18 
  input [18:0] Wgt_4_731, // sfix19_En18 
  input [18:0] Wgt_4_732, // sfix19_En18 
  input [18:0] Wgt_4_733, // sfix19_En18 
  input [18:0] Wgt_4_734, // sfix19_En18 
  input [18:0] Wgt_4_735, // sfix19_En18 
  input [18:0] Wgt_4_736, // sfix19_En18 
  input [18:0] Wgt_4_737, // sfix19_En18 
  input [18:0] Wgt_4_738, // sfix19_En18 
  input [18:0] Wgt_4_739, // sfix19_En18 
  input [18:0] Wgt_4_740, // sfix19_En18 
  input [18:0] Wgt_4_741, // sfix19_En18 
  input [18:0] Wgt_4_742, // sfix19_En18 
  input [18:0] Wgt_4_743, // sfix19_En18 
  input [18:0] Wgt_4_744, // sfix19_En18 
  input [18:0] Wgt_4_745, // sfix19_En18 
  input [18:0] Wgt_4_746, // sfix19_En18 
  input [18:0] Wgt_4_747, // sfix19_En18 
  input [18:0] Wgt_4_748, // sfix19_En18 
  input [18:0] Wgt_4_749, // sfix19_En18 
  input [18:0] Wgt_4_750, // sfix19_En18 
  input [18:0] Wgt_4_751, // sfix19_En18 
  input [18:0] Wgt_4_752, // sfix19_En18 
  input [18:0] Wgt_4_753, // sfix19_En18 
  input [18:0] Wgt_4_754, // sfix19_En18 
  input [18:0] Wgt_4_755, // sfix19_En18 
  input [18:0] Wgt_4_756, // sfix19_En18 
  input [18:0] Wgt_4_757, // sfix19_En18 
  input [18:0] Wgt_4_758, // sfix19_En18 
  input [18:0] Wgt_4_759, // sfix19_En18 
  input [18:0] Wgt_4_760, // sfix19_En18 
  input [18:0] Wgt_4_761, // sfix19_En18 
  input [18:0] Wgt_4_762, // sfix19_En18 
  input [18:0] Wgt_4_763, // sfix19_En18 
  input [18:0] Wgt_4_764, // sfix19_En18 
  input [18:0] Wgt_4_765, // sfix19_En18 
  input [18:0] Wgt_4_766, // sfix19_En18 
  input [18:0] Wgt_4_767, // sfix19_En18 
  input [18:0] Wgt_4_768, // sfix19_En18 
  input [18:0] Wgt_4_769, // sfix19_En18 
  input [18:0] Wgt_4_770, // sfix19_En18 
  input [18:0] Wgt_4_771, // sfix19_En18 
  input [18:0] Wgt_4_772, // sfix19_En18 
  input [18:0] Wgt_4_773, // sfix19_En18 
  input [18:0] Wgt_4_774, // sfix19_En18 
  input [18:0] Wgt_4_775, // sfix19_En18 
  input [18:0] Wgt_4_776, // sfix19_En18 
  input [18:0] Wgt_4_777, // sfix19_En18 
  input [18:0] Wgt_4_778, // sfix19_En18 
  input [18:0] Wgt_4_779, // sfix19_En18 
  input [18:0] Wgt_4_780, // sfix19_En18 
  input [18:0] Wgt_4_781, // sfix19_En18 
  input [18:0] Wgt_4_782, // sfix19_En18 
  input [18:0] Wgt_4_783, // sfix19_En18 
  input [18:0] Wgt_4_784, // sfix19_En18 
  input [18:0] Wgt_5_0, // sfix19_En18 
  input [18:0] Wgt_5_1, // sfix19_En18 
  input [18:0] Wgt_5_2, // sfix19_En18 
  input [18:0] Wgt_5_3, // sfix19_En18 
  input [18:0] Wgt_5_4, // sfix19_En18 
  input [18:0] Wgt_5_5, // sfix19_En18 
  input [18:0] Wgt_5_6, // sfix19_En18 
  input [18:0] Wgt_5_7, // sfix19_En18 
  input [18:0] Wgt_5_8, // sfix19_En18 
  input [18:0] Wgt_5_9, // sfix19_En18 
  input [18:0] Wgt_5_10, // sfix19_En18 
  input [18:0] Wgt_5_11, // sfix19_En18 
  input [18:0] Wgt_5_12, // sfix19_En18 
  input [18:0] Wgt_5_13, // sfix19_En18 
  input [18:0] Wgt_5_14, // sfix19_En18 
  input [18:0] Wgt_5_15, // sfix19_En18 
  input [18:0] Wgt_5_16, // sfix19_En18 
  input [18:0] Wgt_5_17, // sfix19_En18 
  input [18:0] Wgt_5_18, // sfix19_En18 
  input [18:0] Wgt_5_19, // sfix19_En18 
  input [18:0] Wgt_5_20, // sfix19_En18 
  input [18:0] Wgt_5_21, // sfix19_En18 
  input [18:0] Wgt_5_22, // sfix19_En18 
  input [18:0] Wgt_5_23, // sfix19_En18 
  input [18:0] Wgt_5_24, // sfix19_En18 
  input [18:0] Wgt_5_25, // sfix19_En18 
  input [18:0] Wgt_5_26, // sfix19_En18 
  input [18:0] Wgt_5_27, // sfix19_En18 
  input [18:0] Wgt_5_28, // sfix19_En18 
  input [18:0] Wgt_5_29, // sfix19_En18 
  input [18:0] Wgt_5_30, // sfix19_En18 
  input [18:0] Wgt_5_31, // sfix19_En18 
  input [18:0] Wgt_5_32, // sfix19_En18 
  input [18:0] Wgt_5_33, // sfix19_En18 
  input [18:0] Wgt_5_34, // sfix19_En18 
  input [18:0] Wgt_5_35, // sfix19_En18 
  input [18:0] Wgt_5_36, // sfix19_En18 
  input [18:0] Wgt_5_37, // sfix19_En18 
  input [18:0] Wgt_5_38, // sfix19_En18 
  input [18:0] Wgt_5_39, // sfix19_En18 
  input [18:0] Wgt_5_40, // sfix19_En18 
  input [18:0] Wgt_5_41, // sfix19_En18 
  input [18:0] Wgt_5_42, // sfix19_En18 
  input [18:0] Wgt_5_43, // sfix19_En18 
  input [18:0] Wgt_5_44, // sfix19_En18 
  input [18:0] Wgt_5_45, // sfix19_En18 
  input [18:0] Wgt_5_46, // sfix19_En18 
  input [18:0] Wgt_5_47, // sfix19_En18 
  input [18:0] Wgt_5_48, // sfix19_En18 
  input [18:0] Wgt_5_49, // sfix19_En18 
  input [18:0] Wgt_5_50, // sfix19_En18 
  input [18:0] Wgt_5_51, // sfix19_En18 
  input [18:0] Wgt_5_52, // sfix19_En18 
  input [18:0] Wgt_5_53, // sfix19_En18 
  input [18:0] Wgt_5_54, // sfix19_En18 
  input [18:0] Wgt_5_55, // sfix19_En18 
  input [18:0] Wgt_5_56, // sfix19_En18 
  input [18:0] Wgt_5_57, // sfix19_En18 
  input [18:0] Wgt_5_58, // sfix19_En18 
  input [18:0] Wgt_5_59, // sfix19_En18 
  input [18:0] Wgt_5_60, // sfix19_En18 
  input [18:0] Wgt_5_61, // sfix19_En18 
  input [18:0] Wgt_5_62, // sfix19_En18 
  input [18:0] Wgt_5_63, // sfix19_En18 
  input [18:0] Wgt_5_64, // sfix19_En18 
  input [18:0] Wgt_5_65, // sfix19_En18 
  input [18:0] Wgt_5_66, // sfix19_En18 
  input [18:0] Wgt_5_67, // sfix19_En18 
  input [18:0] Wgt_5_68, // sfix19_En18 
  input [18:0] Wgt_5_69, // sfix19_En18 
  input [18:0] Wgt_5_70, // sfix19_En18 
  input [18:0] Wgt_5_71, // sfix19_En18 
  input [18:0] Wgt_5_72, // sfix19_En18 
  input [18:0] Wgt_5_73, // sfix19_En18 
  input [18:0] Wgt_5_74, // sfix19_En18 
  input [18:0] Wgt_5_75, // sfix19_En18 
  input [18:0] Wgt_5_76, // sfix19_En18 
  input [18:0] Wgt_5_77, // sfix19_En18 
  input [18:0] Wgt_5_78, // sfix19_En18 
  input [18:0] Wgt_5_79, // sfix19_En18 
  input [18:0] Wgt_5_80, // sfix19_En18 
  input [18:0] Wgt_5_81, // sfix19_En18 
  input [18:0] Wgt_5_82, // sfix19_En18 
  input [18:0] Wgt_5_83, // sfix19_En18 
  input [18:0] Wgt_5_84, // sfix19_En18 
  input [18:0] Wgt_5_85, // sfix19_En18 
  input [18:0] Wgt_5_86, // sfix19_En18 
  input [18:0] Wgt_5_87, // sfix19_En18 
  input [18:0] Wgt_5_88, // sfix19_En18 
  input [18:0] Wgt_5_89, // sfix19_En18 
  input [18:0] Wgt_5_90, // sfix19_En18 
  input [18:0] Wgt_5_91, // sfix19_En18 
  input [18:0] Wgt_5_92, // sfix19_En18 
  input [18:0] Wgt_5_93, // sfix19_En18 
  input [18:0] Wgt_5_94, // sfix19_En18 
  input [18:0] Wgt_5_95, // sfix19_En18 
  input [18:0] Wgt_5_96, // sfix19_En18 
  input [18:0] Wgt_5_97, // sfix19_En18 
  input [18:0] Wgt_5_98, // sfix19_En18 
  input [18:0] Wgt_5_99, // sfix19_En18 
  input [18:0] Wgt_5_100, // sfix19_En18 
  input [18:0] Wgt_5_101, // sfix19_En18 
  input [18:0] Wgt_5_102, // sfix19_En18 
  input [18:0] Wgt_5_103, // sfix19_En18 
  input [18:0] Wgt_5_104, // sfix19_En18 
  input [18:0] Wgt_5_105, // sfix19_En18 
  input [18:0] Wgt_5_106, // sfix19_En18 
  input [18:0] Wgt_5_107, // sfix19_En18 
  input [18:0] Wgt_5_108, // sfix19_En18 
  input [18:0] Wgt_5_109, // sfix19_En18 
  input [18:0] Wgt_5_110, // sfix19_En18 
  input [18:0] Wgt_5_111, // sfix19_En18 
  input [18:0] Wgt_5_112, // sfix19_En18 
  input [18:0] Wgt_5_113, // sfix19_En18 
  input [18:0] Wgt_5_114, // sfix19_En18 
  input [18:0] Wgt_5_115, // sfix19_En18 
  input [18:0] Wgt_5_116, // sfix19_En18 
  input [18:0] Wgt_5_117, // sfix19_En18 
  input [18:0] Wgt_5_118, // sfix19_En18 
  input [18:0] Wgt_5_119, // sfix19_En18 
  input [18:0] Wgt_5_120, // sfix19_En18 
  input [18:0] Wgt_5_121, // sfix19_En18 
  input [18:0] Wgt_5_122, // sfix19_En18 
  input [18:0] Wgt_5_123, // sfix19_En18 
  input [18:0] Wgt_5_124, // sfix19_En18 
  input [18:0] Wgt_5_125, // sfix19_En18 
  input [18:0] Wgt_5_126, // sfix19_En18 
  input [18:0] Wgt_5_127, // sfix19_En18 
  input [18:0] Wgt_5_128, // sfix19_En18 
  input [18:0] Wgt_5_129, // sfix19_En18 
  input [18:0] Wgt_5_130, // sfix19_En18 
  input [18:0] Wgt_5_131, // sfix19_En18 
  input [18:0] Wgt_5_132, // sfix19_En18 
  input [18:0] Wgt_5_133, // sfix19_En18 
  input [18:0] Wgt_5_134, // sfix19_En18 
  input [18:0] Wgt_5_135, // sfix19_En18 
  input [18:0] Wgt_5_136, // sfix19_En18 
  input [18:0] Wgt_5_137, // sfix19_En18 
  input [18:0] Wgt_5_138, // sfix19_En18 
  input [18:0] Wgt_5_139, // sfix19_En18 
  input [18:0] Wgt_5_140, // sfix19_En18 
  input [18:0] Wgt_5_141, // sfix19_En18 
  input [18:0] Wgt_5_142, // sfix19_En18 
  input [18:0] Wgt_5_143, // sfix19_En18 
  input [18:0] Wgt_5_144, // sfix19_En18 
  input [18:0] Wgt_5_145, // sfix19_En18 
  input [18:0] Wgt_5_146, // sfix19_En18 
  input [18:0] Wgt_5_147, // sfix19_En18 
  input [18:0] Wgt_5_148, // sfix19_En18 
  input [18:0] Wgt_5_149, // sfix19_En18 
  input [18:0] Wgt_5_150, // sfix19_En18 
  input [18:0] Wgt_5_151, // sfix19_En18 
  input [18:0] Wgt_5_152, // sfix19_En18 
  input [18:0] Wgt_5_153, // sfix19_En18 
  input [18:0] Wgt_5_154, // sfix19_En18 
  input [18:0] Wgt_5_155, // sfix19_En18 
  input [18:0] Wgt_5_156, // sfix19_En18 
  input [18:0] Wgt_5_157, // sfix19_En18 
  input [18:0] Wgt_5_158, // sfix19_En18 
  input [18:0] Wgt_5_159, // sfix19_En18 
  input [18:0] Wgt_5_160, // sfix19_En18 
  input [18:0] Wgt_5_161, // sfix19_En18 
  input [18:0] Wgt_5_162, // sfix19_En18 
  input [18:0] Wgt_5_163, // sfix19_En18 
  input [18:0] Wgt_5_164, // sfix19_En18 
  input [18:0] Wgt_5_165, // sfix19_En18 
  input [18:0] Wgt_5_166, // sfix19_En18 
  input [18:0] Wgt_5_167, // sfix19_En18 
  input [18:0] Wgt_5_168, // sfix19_En18 
  input [18:0] Wgt_5_169, // sfix19_En18 
  input [18:0] Wgt_5_170, // sfix19_En18 
  input [18:0] Wgt_5_171, // sfix19_En18 
  input [18:0] Wgt_5_172, // sfix19_En18 
  input [18:0] Wgt_5_173, // sfix19_En18 
  input [18:0] Wgt_5_174, // sfix19_En18 
  input [18:0] Wgt_5_175, // sfix19_En18 
  input [18:0] Wgt_5_176, // sfix19_En18 
  input [18:0] Wgt_5_177, // sfix19_En18 
  input [18:0] Wgt_5_178, // sfix19_En18 
  input [18:0] Wgt_5_179, // sfix19_En18 
  input [18:0] Wgt_5_180, // sfix19_En18 
  input [18:0] Wgt_5_181, // sfix19_En18 
  input [18:0] Wgt_5_182, // sfix19_En18 
  input [18:0] Wgt_5_183, // sfix19_En18 
  input [18:0] Wgt_5_184, // sfix19_En18 
  input [18:0] Wgt_5_185, // sfix19_En18 
  input [18:0] Wgt_5_186, // sfix19_En18 
  input [18:0] Wgt_5_187, // sfix19_En18 
  input [18:0] Wgt_5_188, // sfix19_En18 
  input [18:0] Wgt_5_189, // sfix19_En18 
  input [18:0] Wgt_5_190, // sfix19_En18 
  input [18:0] Wgt_5_191, // sfix19_En18 
  input [18:0] Wgt_5_192, // sfix19_En18 
  input [18:0] Wgt_5_193, // sfix19_En18 
  input [18:0] Wgt_5_194, // sfix19_En18 
  input [18:0] Wgt_5_195, // sfix19_En18 
  input [18:0] Wgt_5_196, // sfix19_En18 
  input [18:0] Wgt_5_197, // sfix19_En18 
  input [18:0] Wgt_5_198, // sfix19_En18 
  input [18:0] Wgt_5_199, // sfix19_En18 
  input [18:0] Wgt_5_200, // sfix19_En18 
  input [18:0] Wgt_5_201, // sfix19_En18 
  input [18:0] Wgt_5_202, // sfix19_En18 
  input [18:0] Wgt_5_203, // sfix19_En18 
  input [18:0] Wgt_5_204, // sfix19_En18 
  input [18:0] Wgt_5_205, // sfix19_En18 
  input [18:0] Wgt_5_206, // sfix19_En18 
  input [18:0] Wgt_5_207, // sfix19_En18 
  input [18:0] Wgt_5_208, // sfix19_En18 
  input [18:0] Wgt_5_209, // sfix19_En18 
  input [18:0] Wgt_5_210, // sfix19_En18 
  input [18:0] Wgt_5_211, // sfix19_En18 
  input [18:0] Wgt_5_212, // sfix19_En18 
  input [18:0] Wgt_5_213, // sfix19_En18 
  input [18:0] Wgt_5_214, // sfix19_En18 
  input [18:0] Wgt_5_215, // sfix19_En18 
  input [18:0] Wgt_5_216, // sfix19_En18 
  input [18:0] Wgt_5_217, // sfix19_En18 
  input [18:0] Wgt_5_218, // sfix19_En18 
  input [18:0] Wgt_5_219, // sfix19_En18 
  input [18:0] Wgt_5_220, // sfix19_En18 
  input [18:0] Wgt_5_221, // sfix19_En18 
  input [18:0] Wgt_5_222, // sfix19_En18 
  input [18:0] Wgt_5_223, // sfix19_En18 
  input [18:0] Wgt_5_224, // sfix19_En18 
  input [18:0] Wgt_5_225, // sfix19_En18 
  input [18:0] Wgt_5_226, // sfix19_En18 
  input [18:0] Wgt_5_227, // sfix19_En18 
  input [18:0] Wgt_5_228, // sfix19_En18 
  input [18:0] Wgt_5_229, // sfix19_En18 
  input [18:0] Wgt_5_230, // sfix19_En18 
  input [18:0] Wgt_5_231, // sfix19_En18 
  input [18:0] Wgt_5_232, // sfix19_En18 
  input [18:0] Wgt_5_233, // sfix19_En18 
  input [18:0] Wgt_5_234, // sfix19_En18 
  input [18:0] Wgt_5_235, // sfix19_En18 
  input [18:0] Wgt_5_236, // sfix19_En18 
  input [18:0] Wgt_5_237, // sfix19_En18 
  input [18:0] Wgt_5_238, // sfix19_En18 
  input [18:0] Wgt_5_239, // sfix19_En18 
  input [18:0] Wgt_5_240, // sfix19_En18 
  input [18:0] Wgt_5_241, // sfix19_En18 
  input [18:0] Wgt_5_242, // sfix19_En18 
  input [18:0] Wgt_5_243, // sfix19_En18 
  input [18:0] Wgt_5_244, // sfix19_En18 
  input [18:0] Wgt_5_245, // sfix19_En18 
  input [18:0] Wgt_5_246, // sfix19_En18 
  input [18:0] Wgt_5_247, // sfix19_En18 
  input [18:0] Wgt_5_248, // sfix19_En18 
  input [18:0] Wgt_5_249, // sfix19_En18 
  input [18:0] Wgt_5_250, // sfix19_En18 
  input [18:0] Wgt_5_251, // sfix19_En18 
  input [18:0] Wgt_5_252, // sfix19_En18 
  input [18:0] Wgt_5_253, // sfix19_En18 
  input [18:0] Wgt_5_254, // sfix19_En18 
  input [18:0] Wgt_5_255, // sfix19_En18 
  input [18:0] Wgt_5_256, // sfix19_En18 
  input [18:0] Wgt_5_257, // sfix19_En18 
  input [18:0] Wgt_5_258, // sfix19_En18 
  input [18:0] Wgt_5_259, // sfix19_En18 
  input [18:0] Wgt_5_260, // sfix19_En18 
  input [18:0] Wgt_5_261, // sfix19_En18 
  input [18:0] Wgt_5_262, // sfix19_En18 
  input [18:0] Wgt_5_263, // sfix19_En18 
  input [18:0] Wgt_5_264, // sfix19_En18 
  input [18:0] Wgt_5_265, // sfix19_En18 
  input [18:0] Wgt_5_266, // sfix19_En18 
  input [18:0] Wgt_5_267, // sfix19_En18 
  input [18:0] Wgt_5_268, // sfix19_En18 
  input [18:0] Wgt_5_269, // sfix19_En18 
  input [18:0] Wgt_5_270, // sfix19_En18 
  input [18:0] Wgt_5_271, // sfix19_En18 
  input [18:0] Wgt_5_272, // sfix19_En18 
  input [18:0] Wgt_5_273, // sfix19_En18 
  input [18:0] Wgt_5_274, // sfix19_En18 
  input [18:0] Wgt_5_275, // sfix19_En18 
  input [18:0] Wgt_5_276, // sfix19_En18 
  input [18:0] Wgt_5_277, // sfix19_En18 
  input [18:0] Wgt_5_278, // sfix19_En18 
  input [18:0] Wgt_5_279, // sfix19_En18 
  input [18:0] Wgt_5_280, // sfix19_En18 
  input [18:0] Wgt_5_281, // sfix19_En18 
  input [18:0] Wgt_5_282, // sfix19_En18 
  input [18:0] Wgt_5_283, // sfix19_En18 
  input [18:0] Wgt_5_284, // sfix19_En18 
  input [18:0] Wgt_5_285, // sfix19_En18 
  input [18:0] Wgt_5_286, // sfix19_En18 
  input [18:0] Wgt_5_287, // sfix19_En18 
  input [18:0] Wgt_5_288, // sfix19_En18 
  input [18:0] Wgt_5_289, // sfix19_En18 
  input [18:0] Wgt_5_290, // sfix19_En18 
  input [18:0] Wgt_5_291, // sfix19_En18 
  input [18:0] Wgt_5_292, // sfix19_En18 
  input [18:0] Wgt_5_293, // sfix19_En18 
  input [18:0] Wgt_5_294, // sfix19_En18 
  input [18:0] Wgt_5_295, // sfix19_En18 
  input [18:0] Wgt_5_296, // sfix19_En18 
  input [18:0] Wgt_5_297, // sfix19_En18 
  input [18:0] Wgt_5_298, // sfix19_En18 
  input [18:0] Wgt_5_299, // sfix19_En18 
  input [18:0] Wgt_5_300, // sfix19_En18 
  input [18:0] Wgt_5_301, // sfix19_En18 
  input [18:0] Wgt_5_302, // sfix19_En18 
  input [18:0] Wgt_5_303, // sfix19_En18 
  input [18:0] Wgt_5_304, // sfix19_En18 
  input [18:0] Wgt_5_305, // sfix19_En18 
  input [18:0] Wgt_5_306, // sfix19_En18 
  input [18:0] Wgt_5_307, // sfix19_En18 
  input [18:0] Wgt_5_308, // sfix19_En18 
  input [18:0] Wgt_5_309, // sfix19_En18 
  input [18:0] Wgt_5_310, // sfix19_En18 
  input [18:0] Wgt_5_311, // sfix19_En18 
  input [18:0] Wgt_5_312, // sfix19_En18 
  input [18:0] Wgt_5_313, // sfix19_En18 
  input [18:0] Wgt_5_314, // sfix19_En18 
  input [18:0] Wgt_5_315, // sfix19_En18 
  input [18:0] Wgt_5_316, // sfix19_En18 
  input [18:0] Wgt_5_317, // sfix19_En18 
  input [18:0] Wgt_5_318, // sfix19_En18 
  input [18:0] Wgt_5_319, // sfix19_En18 
  input [18:0] Wgt_5_320, // sfix19_En18 
  input [18:0] Wgt_5_321, // sfix19_En18 
  input [18:0] Wgt_5_322, // sfix19_En18 
  input [18:0] Wgt_5_323, // sfix19_En18 
  input [18:0] Wgt_5_324, // sfix19_En18 
  input [18:0] Wgt_5_325, // sfix19_En18 
  input [18:0] Wgt_5_326, // sfix19_En18 
  input [18:0] Wgt_5_327, // sfix19_En18 
  input [18:0] Wgt_5_328, // sfix19_En18 
  input [18:0] Wgt_5_329, // sfix19_En18 
  input [18:0] Wgt_5_330, // sfix19_En18 
  input [18:0] Wgt_5_331, // sfix19_En18 
  input [18:0] Wgt_5_332, // sfix19_En18 
  input [18:0] Wgt_5_333, // sfix19_En18 
  input [18:0] Wgt_5_334, // sfix19_En18 
  input [18:0] Wgt_5_335, // sfix19_En18 
  input [18:0] Wgt_5_336, // sfix19_En18 
  input [18:0] Wgt_5_337, // sfix19_En18 
  input [18:0] Wgt_5_338, // sfix19_En18 
  input [18:0] Wgt_5_339, // sfix19_En18 
  input [18:0] Wgt_5_340, // sfix19_En18 
  input [18:0] Wgt_5_341, // sfix19_En18 
  input [18:0] Wgt_5_342, // sfix19_En18 
  input [18:0] Wgt_5_343, // sfix19_En18 
  input [18:0] Wgt_5_344, // sfix19_En18 
  input [18:0] Wgt_5_345, // sfix19_En18 
  input [18:0] Wgt_5_346, // sfix19_En18 
  input [18:0] Wgt_5_347, // sfix19_En18 
  input [18:0] Wgt_5_348, // sfix19_En18 
  input [18:0] Wgt_5_349, // sfix19_En18 
  input [18:0] Wgt_5_350, // sfix19_En18 
  input [18:0] Wgt_5_351, // sfix19_En18 
  input [18:0] Wgt_5_352, // sfix19_En18 
  input [18:0] Wgt_5_353, // sfix19_En18 
  input [18:0] Wgt_5_354, // sfix19_En18 
  input [18:0] Wgt_5_355, // sfix19_En18 
  input [18:0] Wgt_5_356, // sfix19_En18 
  input [18:0] Wgt_5_357, // sfix19_En18 
  input [18:0] Wgt_5_358, // sfix19_En18 
  input [18:0] Wgt_5_359, // sfix19_En18 
  input [18:0] Wgt_5_360, // sfix19_En18 
  input [18:0] Wgt_5_361, // sfix19_En18 
  input [18:0] Wgt_5_362, // sfix19_En18 
  input [18:0] Wgt_5_363, // sfix19_En18 
  input [18:0] Wgt_5_364, // sfix19_En18 
  input [18:0] Wgt_5_365, // sfix19_En18 
  input [18:0] Wgt_5_366, // sfix19_En18 
  input [18:0] Wgt_5_367, // sfix19_En18 
  input [18:0] Wgt_5_368, // sfix19_En18 
  input [18:0] Wgt_5_369, // sfix19_En18 
  input [18:0] Wgt_5_370, // sfix19_En18 
  input [18:0] Wgt_5_371, // sfix19_En18 
  input [18:0] Wgt_5_372, // sfix19_En18 
  input [18:0] Wgt_5_373, // sfix19_En18 
  input [18:0] Wgt_5_374, // sfix19_En18 
  input [18:0] Wgt_5_375, // sfix19_En18 
  input [18:0] Wgt_5_376, // sfix19_En18 
  input [18:0] Wgt_5_377, // sfix19_En18 
  input [18:0] Wgt_5_378, // sfix19_En18 
  input [18:0] Wgt_5_379, // sfix19_En18 
  input [18:0] Wgt_5_380, // sfix19_En18 
  input [18:0] Wgt_5_381, // sfix19_En18 
  input [18:0] Wgt_5_382, // sfix19_En18 
  input [18:0] Wgt_5_383, // sfix19_En18 
  input [18:0] Wgt_5_384, // sfix19_En18 
  input [18:0] Wgt_5_385, // sfix19_En18 
  input [18:0] Wgt_5_386, // sfix19_En18 
  input [18:0] Wgt_5_387, // sfix19_En18 
  input [18:0] Wgt_5_388, // sfix19_En18 
  input [18:0] Wgt_5_389, // sfix19_En18 
  input [18:0] Wgt_5_390, // sfix19_En18 
  input [18:0] Wgt_5_391, // sfix19_En18 
  input [18:0] Wgt_5_392, // sfix19_En18 
  input [18:0] Wgt_5_393, // sfix19_En18 
  input [18:0] Wgt_5_394, // sfix19_En18 
  input [18:0] Wgt_5_395, // sfix19_En18 
  input [18:0] Wgt_5_396, // sfix19_En18 
  input [18:0] Wgt_5_397, // sfix19_En18 
  input [18:0] Wgt_5_398, // sfix19_En18 
  input [18:0] Wgt_5_399, // sfix19_En18 
  input [18:0] Wgt_5_400, // sfix19_En18 
  input [18:0] Wgt_5_401, // sfix19_En18 
  input [18:0] Wgt_5_402, // sfix19_En18 
  input [18:0] Wgt_5_403, // sfix19_En18 
  input [18:0] Wgt_5_404, // sfix19_En18 
  input [18:0] Wgt_5_405, // sfix19_En18 
  input [18:0] Wgt_5_406, // sfix19_En18 
  input [18:0] Wgt_5_407, // sfix19_En18 
  input [18:0] Wgt_5_408, // sfix19_En18 
  input [18:0] Wgt_5_409, // sfix19_En18 
  input [18:0] Wgt_5_410, // sfix19_En18 
  input [18:0] Wgt_5_411, // sfix19_En18 
  input [18:0] Wgt_5_412, // sfix19_En18 
  input [18:0] Wgt_5_413, // sfix19_En18 
  input [18:0] Wgt_5_414, // sfix19_En18 
  input [18:0] Wgt_5_415, // sfix19_En18 
  input [18:0] Wgt_5_416, // sfix19_En18 
  input [18:0] Wgt_5_417, // sfix19_En18 
  input [18:0] Wgt_5_418, // sfix19_En18 
  input [18:0] Wgt_5_419, // sfix19_En18 
  input [18:0] Wgt_5_420, // sfix19_En18 
  input [18:0] Wgt_5_421, // sfix19_En18 
  input [18:0] Wgt_5_422, // sfix19_En18 
  input [18:0] Wgt_5_423, // sfix19_En18 
  input [18:0] Wgt_5_424, // sfix19_En18 
  input [18:0] Wgt_5_425, // sfix19_En18 
  input [18:0] Wgt_5_426, // sfix19_En18 
  input [18:0] Wgt_5_427, // sfix19_En18 
  input [18:0] Wgt_5_428, // sfix19_En18 
  input [18:0] Wgt_5_429, // sfix19_En18 
  input [18:0] Wgt_5_430, // sfix19_En18 
  input [18:0] Wgt_5_431, // sfix19_En18 
  input [18:0] Wgt_5_432, // sfix19_En18 
  input [18:0] Wgt_5_433, // sfix19_En18 
  input [18:0] Wgt_5_434, // sfix19_En18 
  input [18:0] Wgt_5_435, // sfix19_En18 
  input [18:0] Wgt_5_436, // sfix19_En18 
  input [18:0] Wgt_5_437, // sfix19_En18 
  input [18:0] Wgt_5_438, // sfix19_En18 
  input [18:0] Wgt_5_439, // sfix19_En18 
  input [18:0] Wgt_5_440, // sfix19_En18 
  input [18:0] Wgt_5_441, // sfix19_En18 
  input [18:0] Wgt_5_442, // sfix19_En18 
  input [18:0] Wgt_5_443, // sfix19_En18 
  input [18:0] Wgt_5_444, // sfix19_En18 
  input [18:0] Wgt_5_445, // sfix19_En18 
  input [18:0] Wgt_5_446, // sfix19_En18 
  input [18:0] Wgt_5_447, // sfix19_En18 
  input [18:0] Wgt_5_448, // sfix19_En18 
  input [18:0] Wgt_5_449, // sfix19_En18 
  input [18:0] Wgt_5_450, // sfix19_En18 
  input [18:0] Wgt_5_451, // sfix19_En18 
  input [18:0] Wgt_5_452, // sfix19_En18 
  input [18:0] Wgt_5_453, // sfix19_En18 
  input [18:0] Wgt_5_454, // sfix19_En18 
  input [18:0] Wgt_5_455, // sfix19_En18 
  input [18:0] Wgt_5_456, // sfix19_En18 
  input [18:0] Wgt_5_457, // sfix19_En18 
  input [18:0] Wgt_5_458, // sfix19_En18 
  input [18:0] Wgt_5_459, // sfix19_En18 
  input [18:0] Wgt_5_460, // sfix19_En18 
  input [18:0] Wgt_5_461, // sfix19_En18 
  input [18:0] Wgt_5_462, // sfix19_En18 
  input [18:0] Wgt_5_463, // sfix19_En18 
  input [18:0] Wgt_5_464, // sfix19_En18 
  input [18:0] Wgt_5_465, // sfix19_En18 
  input [18:0] Wgt_5_466, // sfix19_En18 
  input [18:0] Wgt_5_467, // sfix19_En18 
  input [18:0] Wgt_5_468, // sfix19_En18 
  input [18:0] Wgt_5_469, // sfix19_En18 
  input [18:0] Wgt_5_470, // sfix19_En18 
  input [18:0] Wgt_5_471, // sfix19_En18 
  input [18:0] Wgt_5_472, // sfix19_En18 
  input [18:0] Wgt_5_473, // sfix19_En18 
  input [18:0] Wgt_5_474, // sfix19_En18 
  input [18:0] Wgt_5_475, // sfix19_En18 
  input [18:0] Wgt_5_476, // sfix19_En18 
  input [18:0] Wgt_5_477, // sfix19_En18 
  input [18:0] Wgt_5_478, // sfix19_En18 
  input [18:0] Wgt_5_479, // sfix19_En18 
  input [18:0] Wgt_5_480, // sfix19_En18 
  input [18:0] Wgt_5_481, // sfix19_En18 
  input [18:0] Wgt_5_482, // sfix19_En18 
  input [18:0] Wgt_5_483, // sfix19_En18 
  input [18:0] Wgt_5_484, // sfix19_En18 
  input [18:0] Wgt_5_485, // sfix19_En18 
  input [18:0] Wgt_5_486, // sfix19_En18 
  input [18:0] Wgt_5_487, // sfix19_En18 
  input [18:0] Wgt_5_488, // sfix19_En18 
  input [18:0] Wgt_5_489, // sfix19_En18 
  input [18:0] Wgt_5_490, // sfix19_En18 
  input [18:0] Wgt_5_491, // sfix19_En18 
  input [18:0] Wgt_5_492, // sfix19_En18 
  input [18:0] Wgt_5_493, // sfix19_En18 
  input [18:0] Wgt_5_494, // sfix19_En18 
  input [18:0] Wgt_5_495, // sfix19_En18 
  input [18:0] Wgt_5_496, // sfix19_En18 
  input [18:0] Wgt_5_497, // sfix19_En18 
  input [18:0] Wgt_5_498, // sfix19_En18 
  input [18:0] Wgt_5_499, // sfix19_En18 
  input [18:0] Wgt_5_500, // sfix19_En18 
  input [18:0] Wgt_5_501, // sfix19_En18 
  input [18:0] Wgt_5_502, // sfix19_En18 
  input [18:0] Wgt_5_503, // sfix19_En18 
  input [18:0] Wgt_5_504, // sfix19_En18 
  input [18:0] Wgt_5_505, // sfix19_En18 
  input [18:0] Wgt_5_506, // sfix19_En18 
  input [18:0] Wgt_5_507, // sfix19_En18 
  input [18:0] Wgt_5_508, // sfix19_En18 
  input [18:0] Wgt_5_509, // sfix19_En18 
  input [18:0] Wgt_5_510, // sfix19_En18 
  input [18:0] Wgt_5_511, // sfix19_En18 
  input [18:0] Wgt_5_512, // sfix19_En18 
  input [18:0] Wgt_5_513, // sfix19_En18 
  input [18:0] Wgt_5_514, // sfix19_En18 
  input [18:0] Wgt_5_515, // sfix19_En18 
  input [18:0] Wgt_5_516, // sfix19_En18 
  input [18:0] Wgt_5_517, // sfix19_En18 
  input [18:0] Wgt_5_518, // sfix19_En18 
  input [18:0] Wgt_5_519, // sfix19_En18 
  input [18:0] Wgt_5_520, // sfix19_En18 
  input [18:0] Wgt_5_521, // sfix19_En18 
  input [18:0] Wgt_5_522, // sfix19_En18 
  input [18:0] Wgt_5_523, // sfix19_En18 
  input [18:0] Wgt_5_524, // sfix19_En18 
  input [18:0] Wgt_5_525, // sfix19_En18 
  input [18:0] Wgt_5_526, // sfix19_En18 
  input [18:0] Wgt_5_527, // sfix19_En18 
  input [18:0] Wgt_5_528, // sfix19_En18 
  input [18:0] Wgt_5_529, // sfix19_En18 
  input [18:0] Wgt_5_530, // sfix19_En18 
  input [18:0] Wgt_5_531, // sfix19_En18 
  input [18:0] Wgt_5_532, // sfix19_En18 
  input [18:0] Wgt_5_533, // sfix19_En18 
  input [18:0] Wgt_5_534, // sfix19_En18 
  input [18:0] Wgt_5_535, // sfix19_En18 
  input [18:0] Wgt_5_536, // sfix19_En18 
  input [18:0] Wgt_5_537, // sfix19_En18 
  input [18:0] Wgt_5_538, // sfix19_En18 
  input [18:0] Wgt_5_539, // sfix19_En18 
  input [18:0] Wgt_5_540, // sfix19_En18 
  input [18:0] Wgt_5_541, // sfix19_En18 
  input [18:0] Wgt_5_542, // sfix19_En18 
  input [18:0] Wgt_5_543, // sfix19_En18 
  input [18:0] Wgt_5_544, // sfix19_En18 
  input [18:0] Wgt_5_545, // sfix19_En18 
  input [18:0] Wgt_5_546, // sfix19_En18 
  input [18:0] Wgt_5_547, // sfix19_En18 
  input [18:0] Wgt_5_548, // sfix19_En18 
  input [18:0] Wgt_5_549, // sfix19_En18 
  input [18:0] Wgt_5_550, // sfix19_En18 
  input [18:0] Wgt_5_551, // sfix19_En18 
  input [18:0] Wgt_5_552, // sfix19_En18 
  input [18:0] Wgt_5_553, // sfix19_En18 
  input [18:0] Wgt_5_554, // sfix19_En18 
  input [18:0] Wgt_5_555, // sfix19_En18 
  input [18:0] Wgt_5_556, // sfix19_En18 
  input [18:0] Wgt_5_557, // sfix19_En18 
  input [18:0] Wgt_5_558, // sfix19_En18 
  input [18:0] Wgt_5_559, // sfix19_En18 
  input [18:0] Wgt_5_560, // sfix19_En18 
  input [18:0] Wgt_5_561, // sfix19_En18 
  input [18:0] Wgt_5_562, // sfix19_En18 
  input [18:0] Wgt_5_563, // sfix19_En18 
  input [18:0] Wgt_5_564, // sfix19_En18 
  input [18:0] Wgt_5_565, // sfix19_En18 
  input [18:0] Wgt_5_566, // sfix19_En18 
  input [18:0] Wgt_5_567, // sfix19_En18 
  input [18:0] Wgt_5_568, // sfix19_En18 
  input [18:0] Wgt_5_569, // sfix19_En18 
  input [18:0] Wgt_5_570, // sfix19_En18 
  input [18:0] Wgt_5_571, // sfix19_En18 
  input [18:0] Wgt_5_572, // sfix19_En18 
  input [18:0] Wgt_5_573, // sfix19_En18 
  input [18:0] Wgt_5_574, // sfix19_En18 
  input [18:0] Wgt_5_575, // sfix19_En18 
  input [18:0] Wgt_5_576, // sfix19_En18 
  input [18:0] Wgt_5_577, // sfix19_En18 
  input [18:0] Wgt_5_578, // sfix19_En18 
  input [18:0] Wgt_5_579, // sfix19_En18 
  input [18:0] Wgt_5_580, // sfix19_En18 
  input [18:0] Wgt_5_581, // sfix19_En18 
  input [18:0] Wgt_5_582, // sfix19_En18 
  input [18:0] Wgt_5_583, // sfix19_En18 
  input [18:0] Wgt_5_584, // sfix19_En18 
  input [18:0] Wgt_5_585, // sfix19_En18 
  input [18:0] Wgt_5_586, // sfix19_En18 
  input [18:0] Wgt_5_587, // sfix19_En18 
  input [18:0] Wgt_5_588, // sfix19_En18 
  input [18:0] Wgt_5_589, // sfix19_En18 
  input [18:0] Wgt_5_590, // sfix19_En18 
  input [18:0] Wgt_5_591, // sfix19_En18 
  input [18:0] Wgt_5_592, // sfix19_En18 
  input [18:0] Wgt_5_593, // sfix19_En18 
  input [18:0] Wgt_5_594, // sfix19_En18 
  input [18:0] Wgt_5_595, // sfix19_En18 
  input [18:0] Wgt_5_596, // sfix19_En18 
  input [18:0] Wgt_5_597, // sfix19_En18 
  input [18:0] Wgt_5_598, // sfix19_En18 
  input [18:0] Wgt_5_599, // sfix19_En18 
  input [18:0] Wgt_5_600, // sfix19_En18 
  input [18:0] Wgt_5_601, // sfix19_En18 
  input [18:0] Wgt_5_602, // sfix19_En18 
  input [18:0] Wgt_5_603, // sfix19_En18 
  input [18:0] Wgt_5_604, // sfix19_En18 
  input [18:0] Wgt_5_605, // sfix19_En18 
  input [18:0] Wgt_5_606, // sfix19_En18 
  input [18:0] Wgt_5_607, // sfix19_En18 
  input [18:0] Wgt_5_608, // sfix19_En18 
  input [18:0] Wgt_5_609, // sfix19_En18 
  input [18:0] Wgt_5_610, // sfix19_En18 
  input [18:0] Wgt_5_611, // sfix19_En18 
  input [18:0] Wgt_5_612, // sfix19_En18 
  input [18:0] Wgt_5_613, // sfix19_En18 
  input [18:0] Wgt_5_614, // sfix19_En18 
  input [18:0] Wgt_5_615, // sfix19_En18 
  input [18:0] Wgt_5_616, // sfix19_En18 
  input [18:0] Wgt_5_617, // sfix19_En18 
  input [18:0] Wgt_5_618, // sfix19_En18 
  input [18:0] Wgt_5_619, // sfix19_En18 
  input [18:0] Wgt_5_620, // sfix19_En18 
  input [18:0] Wgt_5_621, // sfix19_En18 
  input [18:0] Wgt_5_622, // sfix19_En18 
  input [18:0] Wgt_5_623, // sfix19_En18 
  input [18:0] Wgt_5_624, // sfix19_En18 
  input [18:0] Wgt_5_625, // sfix19_En18 
  input [18:0] Wgt_5_626, // sfix19_En18 
  input [18:0] Wgt_5_627, // sfix19_En18 
  input [18:0] Wgt_5_628, // sfix19_En18 
  input [18:0] Wgt_5_629, // sfix19_En18 
  input [18:0] Wgt_5_630, // sfix19_En18 
  input [18:0] Wgt_5_631, // sfix19_En18 
  input [18:0] Wgt_5_632, // sfix19_En18 
  input [18:0] Wgt_5_633, // sfix19_En18 
  input [18:0] Wgt_5_634, // sfix19_En18 
  input [18:0] Wgt_5_635, // sfix19_En18 
  input [18:0] Wgt_5_636, // sfix19_En18 
  input [18:0] Wgt_5_637, // sfix19_En18 
  input [18:0] Wgt_5_638, // sfix19_En18 
  input [18:0] Wgt_5_639, // sfix19_En18 
  input [18:0] Wgt_5_640, // sfix19_En18 
  input [18:0] Wgt_5_641, // sfix19_En18 
  input [18:0] Wgt_5_642, // sfix19_En18 
  input [18:0] Wgt_5_643, // sfix19_En18 
  input [18:0] Wgt_5_644, // sfix19_En18 
  input [18:0] Wgt_5_645, // sfix19_En18 
  input [18:0] Wgt_5_646, // sfix19_En18 
  input [18:0] Wgt_5_647, // sfix19_En18 
  input [18:0] Wgt_5_648, // sfix19_En18 
  input [18:0] Wgt_5_649, // sfix19_En18 
  input [18:0] Wgt_5_650, // sfix19_En18 
  input [18:0] Wgt_5_651, // sfix19_En18 
  input [18:0] Wgt_5_652, // sfix19_En18 
  input [18:0] Wgt_5_653, // sfix19_En18 
  input [18:0] Wgt_5_654, // sfix19_En18 
  input [18:0] Wgt_5_655, // sfix19_En18 
  input [18:0] Wgt_5_656, // sfix19_En18 
  input [18:0] Wgt_5_657, // sfix19_En18 
  input [18:0] Wgt_5_658, // sfix19_En18 
  input [18:0] Wgt_5_659, // sfix19_En18 
  input [18:0] Wgt_5_660, // sfix19_En18 
  input [18:0] Wgt_5_661, // sfix19_En18 
  input [18:0] Wgt_5_662, // sfix19_En18 
  input [18:0] Wgt_5_663, // sfix19_En18 
  input [18:0] Wgt_5_664, // sfix19_En18 
  input [18:0] Wgt_5_665, // sfix19_En18 
  input [18:0] Wgt_5_666, // sfix19_En18 
  input [18:0] Wgt_5_667, // sfix19_En18 
  input [18:0] Wgt_5_668, // sfix19_En18 
  input [18:0] Wgt_5_669, // sfix19_En18 
  input [18:0] Wgt_5_670, // sfix19_En18 
  input [18:0] Wgt_5_671, // sfix19_En18 
  input [18:0] Wgt_5_672, // sfix19_En18 
  input [18:0] Wgt_5_673, // sfix19_En18 
  input [18:0] Wgt_5_674, // sfix19_En18 
  input [18:0] Wgt_5_675, // sfix19_En18 
  input [18:0] Wgt_5_676, // sfix19_En18 
  input [18:0] Wgt_5_677, // sfix19_En18 
  input [18:0] Wgt_5_678, // sfix19_En18 
  input [18:0] Wgt_5_679, // sfix19_En18 
  input [18:0] Wgt_5_680, // sfix19_En18 
  input [18:0] Wgt_5_681, // sfix19_En18 
  input [18:0] Wgt_5_682, // sfix19_En18 
  input [18:0] Wgt_5_683, // sfix19_En18 
  input [18:0] Wgt_5_684, // sfix19_En18 
  input [18:0] Wgt_5_685, // sfix19_En18 
  input [18:0] Wgt_5_686, // sfix19_En18 
  input [18:0] Wgt_5_687, // sfix19_En18 
  input [18:0] Wgt_5_688, // sfix19_En18 
  input [18:0] Wgt_5_689, // sfix19_En18 
  input [18:0] Wgt_5_690, // sfix19_En18 
  input [18:0] Wgt_5_691, // sfix19_En18 
  input [18:0] Wgt_5_692, // sfix19_En18 
  input [18:0] Wgt_5_693, // sfix19_En18 
  input [18:0] Wgt_5_694, // sfix19_En18 
  input [18:0] Wgt_5_695, // sfix19_En18 
  input [18:0] Wgt_5_696, // sfix19_En18 
  input [18:0] Wgt_5_697, // sfix19_En18 
  input [18:0] Wgt_5_698, // sfix19_En18 
  input [18:0] Wgt_5_699, // sfix19_En18 
  input [18:0] Wgt_5_700, // sfix19_En18 
  input [18:0] Wgt_5_701, // sfix19_En18 
  input [18:0] Wgt_5_702, // sfix19_En18 
  input [18:0] Wgt_5_703, // sfix19_En18 
  input [18:0] Wgt_5_704, // sfix19_En18 
  input [18:0] Wgt_5_705, // sfix19_En18 
  input [18:0] Wgt_5_706, // sfix19_En18 
  input [18:0] Wgt_5_707, // sfix19_En18 
  input [18:0] Wgt_5_708, // sfix19_En18 
  input [18:0] Wgt_5_709, // sfix19_En18 
  input [18:0] Wgt_5_710, // sfix19_En18 
  input [18:0] Wgt_5_711, // sfix19_En18 
  input [18:0] Wgt_5_712, // sfix19_En18 
  input [18:0] Wgt_5_713, // sfix19_En18 
  input [18:0] Wgt_5_714, // sfix19_En18 
  input [18:0] Wgt_5_715, // sfix19_En18 
  input [18:0] Wgt_5_716, // sfix19_En18 
  input [18:0] Wgt_5_717, // sfix19_En18 
  input [18:0] Wgt_5_718, // sfix19_En18 
  input [18:0] Wgt_5_719, // sfix19_En18 
  input [18:0] Wgt_5_720, // sfix19_En18 
  input [18:0] Wgt_5_721, // sfix19_En18 
  input [18:0] Wgt_5_722, // sfix19_En18 
  input [18:0] Wgt_5_723, // sfix19_En18 
  input [18:0] Wgt_5_724, // sfix19_En18 
  input [18:0] Wgt_5_725, // sfix19_En18 
  input [18:0] Wgt_5_726, // sfix19_En18 
  input [18:0] Wgt_5_727, // sfix19_En18 
  input [18:0] Wgt_5_728, // sfix19_En18 
  input [18:0] Wgt_5_729, // sfix19_En18 
  input [18:0] Wgt_5_730, // sfix19_En18 
  input [18:0] Wgt_5_731, // sfix19_En18 
  input [18:0] Wgt_5_732, // sfix19_En18 
  input [18:0] Wgt_5_733, // sfix19_En18 
  input [18:0] Wgt_5_734, // sfix19_En18 
  input [18:0] Wgt_5_735, // sfix19_En18 
  input [18:0] Wgt_5_736, // sfix19_En18 
  input [18:0] Wgt_5_737, // sfix19_En18 
  input [18:0] Wgt_5_738, // sfix19_En18 
  input [18:0] Wgt_5_739, // sfix19_En18 
  input [18:0] Wgt_5_740, // sfix19_En18 
  input [18:0] Wgt_5_741, // sfix19_En18 
  input [18:0] Wgt_5_742, // sfix19_En18 
  input [18:0] Wgt_5_743, // sfix19_En18 
  input [18:0] Wgt_5_744, // sfix19_En18 
  input [18:0] Wgt_5_745, // sfix19_En18 
  input [18:0] Wgt_5_746, // sfix19_En18 
  input [18:0] Wgt_5_747, // sfix19_En18 
  input [18:0] Wgt_5_748, // sfix19_En18 
  input [18:0] Wgt_5_749, // sfix19_En18 
  input [18:0] Wgt_5_750, // sfix19_En18 
  input [18:0] Wgt_5_751, // sfix19_En18 
  input [18:0] Wgt_5_752, // sfix19_En18 
  input [18:0] Wgt_5_753, // sfix19_En18 
  input [18:0] Wgt_5_754, // sfix19_En18 
  input [18:0] Wgt_5_755, // sfix19_En18 
  input [18:0] Wgt_5_756, // sfix19_En18 
  input [18:0] Wgt_5_757, // sfix19_En18 
  input [18:0] Wgt_5_758, // sfix19_En18 
  input [18:0] Wgt_5_759, // sfix19_En18 
  input [18:0] Wgt_5_760, // sfix19_En18 
  input [18:0] Wgt_5_761, // sfix19_En18 
  input [18:0] Wgt_5_762, // sfix19_En18 
  input [18:0] Wgt_5_763, // sfix19_En18 
  input [18:0] Wgt_5_764, // sfix19_En18 
  input [18:0] Wgt_5_765, // sfix19_En18 
  input [18:0] Wgt_5_766, // sfix19_En18 
  input [18:0] Wgt_5_767, // sfix19_En18 
  input [18:0] Wgt_5_768, // sfix19_En18 
  input [18:0] Wgt_5_769, // sfix19_En18 
  input [18:0] Wgt_5_770, // sfix19_En18 
  input [18:0] Wgt_5_771, // sfix19_En18 
  input [18:0] Wgt_5_772, // sfix19_En18 
  input [18:0] Wgt_5_773, // sfix19_En18 
  input [18:0] Wgt_5_774, // sfix19_En18 
  input [18:0] Wgt_5_775, // sfix19_En18 
  input [18:0] Wgt_5_776, // sfix19_En18 
  input [18:0] Wgt_5_777, // sfix19_En18 
  input [18:0] Wgt_5_778, // sfix19_En18 
  input [18:0] Wgt_5_779, // sfix19_En18 
  input [18:0] Wgt_5_780, // sfix19_En18 
  input [18:0] Wgt_5_781, // sfix19_En18 
  input [18:0] Wgt_5_782, // sfix19_En18 
  input [18:0] Wgt_5_783, // sfix19_En18 
  input [18:0] Wgt_5_784, // sfix19_En18 
  input [18:0] Wgt_6_0, // sfix19_En18 
  input [18:0] Wgt_6_1, // sfix19_En18 
  input [18:0] Wgt_6_2, // sfix19_En18 
  input [18:0] Wgt_6_3, // sfix19_En18 
  input [18:0] Wgt_6_4, // sfix19_En18 
  input [18:0] Wgt_6_5, // sfix19_En18 
  input [18:0] Wgt_6_6, // sfix19_En18 
  input [18:0] Wgt_6_7, // sfix19_En18 
  input [18:0] Wgt_6_8, // sfix19_En18 
  input [18:0] Wgt_6_9, // sfix19_En18 
  input [18:0] Wgt_6_10, // sfix19_En18 
  input [18:0] Wgt_6_11, // sfix19_En18 
  input [18:0] Wgt_6_12, // sfix19_En18 
  input [18:0] Wgt_6_13, // sfix19_En18 
  input [18:0] Wgt_6_14, // sfix19_En18 
  input [18:0] Wgt_6_15, // sfix19_En18 
  input [18:0] Wgt_6_16, // sfix19_En18 
  input [18:0] Wgt_6_17, // sfix19_En18 
  input [18:0] Wgt_6_18, // sfix19_En18 
  input [18:0] Wgt_6_19, // sfix19_En18 
  input [18:0] Wgt_6_20, // sfix19_En18 
  input [18:0] Wgt_6_21, // sfix19_En18 
  input [18:0] Wgt_6_22, // sfix19_En18 
  input [18:0] Wgt_6_23, // sfix19_En18 
  input [18:0] Wgt_6_24, // sfix19_En18 
  input [18:0] Wgt_6_25, // sfix19_En18 
  input [18:0] Wgt_6_26, // sfix19_En18 
  input [18:0] Wgt_6_27, // sfix19_En18 
  input [18:0] Wgt_6_28, // sfix19_En18 
  input [18:0] Wgt_6_29, // sfix19_En18 
  input [18:0] Wgt_6_30, // sfix19_En18 
  input [18:0] Wgt_6_31, // sfix19_En18 
  input [18:0] Wgt_6_32, // sfix19_En18 
  input [18:0] Wgt_6_33, // sfix19_En18 
  input [18:0] Wgt_6_34, // sfix19_En18 
  input [18:0] Wgt_6_35, // sfix19_En18 
  input [18:0] Wgt_6_36, // sfix19_En18 
  input [18:0] Wgt_6_37, // sfix19_En18 
  input [18:0] Wgt_6_38, // sfix19_En18 
  input [18:0] Wgt_6_39, // sfix19_En18 
  input [18:0] Wgt_6_40, // sfix19_En18 
  input [18:0] Wgt_6_41, // sfix19_En18 
  input [18:0] Wgt_6_42, // sfix19_En18 
  input [18:0] Wgt_6_43, // sfix19_En18 
  input [18:0] Wgt_6_44, // sfix19_En18 
  input [18:0] Wgt_6_45, // sfix19_En18 
  input [18:0] Wgt_6_46, // sfix19_En18 
  input [18:0] Wgt_6_47, // sfix19_En18 
  input [18:0] Wgt_6_48, // sfix19_En18 
  input [18:0] Wgt_6_49, // sfix19_En18 
  input [18:0] Wgt_6_50, // sfix19_En18 
  input [18:0] Wgt_6_51, // sfix19_En18 
  input [18:0] Wgt_6_52, // sfix19_En18 
  input [18:0] Wgt_6_53, // sfix19_En18 
  input [18:0] Wgt_6_54, // sfix19_En18 
  input [18:0] Wgt_6_55, // sfix19_En18 
  input [18:0] Wgt_6_56, // sfix19_En18 
  input [18:0] Wgt_6_57, // sfix19_En18 
  input [18:0] Wgt_6_58, // sfix19_En18 
  input [18:0] Wgt_6_59, // sfix19_En18 
  input [18:0] Wgt_6_60, // sfix19_En18 
  input [18:0] Wgt_6_61, // sfix19_En18 
  input [18:0] Wgt_6_62, // sfix19_En18 
  input [18:0] Wgt_6_63, // sfix19_En18 
  input [18:0] Wgt_6_64, // sfix19_En18 
  input [18:0] Wgt_6_65, // sfix19_En18 
  input [18:0] Wgt_6_66, // sfix19_En18 
  input [18:0] Wgt_6_67, // sfix19_En18 
  input [18:0] Wgt_6_68, // sfix19_En18 
  input [18:0] Wgt_6_69, // sfix19_En18 
  input [18:0] Wgt_6_70, // sfix19_En18 
  input [18:0] Wgt_6_71, // sfix19_En18 
  input [18:0] Wgt_6_72, // sfix19_En18 
  input [18:0] Wgt_6_73, // sfix19_En18 
  input [18:0] Wgt_6_74, // sfix19_En18 
  input [18:0] Wgt_6_75, // sfix19_En18 
  input [18:0] Wgt_6_76, // sfix19_En18 
  input [18:0] Wgt_6_77, // sfix19_En18 
  input [18:0] Wgt_6_78, // sfix19_En18 
  input [18:0] Wgt_6_79, // sfix19_En18 
  input [18:0] Wgt_6_80, // sfix19_En18 
  input [18:0] Wgt_6_81, // sfix19_En18 
  input [18:0] Wgt_6_82, // sfix19_En18 
  input [18:0] Wgt_6_83, // sfix19_En18 
  input [18:0] Wgt_6_84, // sfix19_En18 
  input [18:0] Wgt_6_85, // sfix19_En18 
  input [18:0] Wgt_6_86, // sfix19_En18 
  input [18:0] Wgt_6_87, // sfix19_En18 
  input [18:0] Wgt_6_88, // sfix19_En18 
  input [18:0] Wgt_6_89, // sfix19_En18 
  input [18:0] Wgt_6_90, // sfix19_En18 
  input [18:0] Wgt_6_91, // sfix19_En18 
  input [18:0] Wgt_6_92, // sfix19_En18 
  input [18:0] Wgt_6_93, // sfix19_En18 
  input [18:0] Wgt_6_94, // sfix19_En18 
  input [18:0] Wgt_6_95, // sfix19_En18 
  input [18:0] Wgt_6_96, // sfix19_En18 
  input [18:0] Wgt_6_97, // sfix19_En18 
  input [18:0] Wgt_6_98, // sfix19_En18 
  input [18:0] Wgt_6_99, // sfix19_En18 
  input [18:0] Wgt_6_100, // sfix19_En18 
  input [18:0] Wgt_6_101, // sfix19_En18 
  input [18:0] Wgt_6_102, // sfix19_En18 
  input [18:0] Wgt_6_103, // sfix19_En18 
  input [18:0] Wgt_6_104, // sfix19_En18 
  input [18:0] Wgt_6_105, // sfix19_En18 
  input [18:0] Wgt_6_106, // sfix19_En18 
  input [18:0] Wgt_6_107, // sfix19_En18 
  input [18:0] Wgt_6_108, // sfix19_En18 
  input [18:0] Wgt_6_109, // sfix19_En18 
  input [18:0] Wgt_6_110, // sfix19_En18 
  input [18:0] Wgt_6_111, // sfix19_En18 
  input [18:0] Wgt_6_112, // sfix19_En18 
  input [18:0] Wgt_6_113, // sfix19_En18 
  input [18:0] Wgt_6_114, // sfix19_En18 
  input [18:0] Wgt_6_115, // sfix19_En18 
  input [18:0] Wgt_6_116, // sfix19_En18 
  input [18:0] Wgt_6_117, // sfix19_En18 
  input [18:0] Wgt_6_118, // sfix19_En18 
  input [18:0] Wgt_6_119, // sfix19_En18 
  input [18:0] Wgt_6_120, // sfix19_En18 
  input [18:0] Wgt_6_121, // sfix19_En18 
  input [18:0] Wgt_6_122, // sfix19_En18 
  input [18:0] Wgt_6_123, // sfix19_En18 
  input [18:0] Wgt_6_124, // sfix19_En18 
  input [18:0] Wgt_6_125, // sfix19_En18 
  input [18:0] Wgt_6_126, // sfix19_En18 
  input [18:0] Wgt_6_127, // sfix19_En18 
  input [18:0] Wgt_6_128, // sfix19_En18 
  input [18:0] Wgt_6_129, // sfix19_En18 
  input [18:0] Wgt_6_130, // sfix19_En18 
  input [18:0] Wgt_6_131, // sfix19_En18 
  input [18:0] Wgt_6_132, // sfix19_En18 
  input [18:0] Wgt_6_133, // sfix19_En18 
  input [18:0] Wgt_6_134, // sfix19_En18 
  input [18:0] Wgt_6_135, // sfix19_En18 
  input [18:0] Wgt_6_136, // sfix19_En18 
  input [18:0] Wgt_6_137, // sfix19_En18 
  input [18:0] Wgt_6_138, // sfix19_En18 
  input [18:0] Wgt_6_139, // sfix19_En18 
  input [18:0] Wgt_6_140, // sfix19_En18 
  input [18:0] Wgt_6_141, // sfix19_En18 
  input [18:0] Wgt_6_142, // sfix19_En18 
  input [18:0] Wgt_6_143, // sfix19_En18 
  input [18:0] Wgt_6_144, // sfix19_En18 
  input [18:0] Wgt_6_145, // sfix19_En18 
  input [18:0] Wgt_6_146, // sfix19_En18 
  input [18:0] Wgt_6_147, // sfix19_En18 
  input [18:0] Wgt_6_148, // sfix19_En18 
  input [18:0] Wgt_6_149, // sfix19_En18 
  input [18:0] Wgt_6_150, // sfix19_En18 
  input [18:0] Wgt_6_151, // sfix19_En18 
  input [18:0] Wgt_6_152, // sfix19_En18 
  input [18:0] Wgt_6_153, // sfix19_En18 
  input [18:0] Wgt_6_154, // sfix19_En18 
  input [18:0] Wgt_6_155, // sfix19_En18 
  input [18:0] Wgt_6_156, // sfix19_En18 
  input [18:0] Wgt_6_157, // sfix19_En18 
  input [18:0] Wgt_6_158, // sfix19_En18 
  input [18:0] Wgt_6_159, // sfix19_En18 
  input [18:0] Wgt_6_160, // sfix19_En18 
  input [18:0] Wgt_6_161, // sfix19_En18 
  input [18:0] Wgt_6_162, // sfix19_En18 
  input [18:0] Wgt_6_163, // sfix19_En18 
  input [18:0] Wgt_6_164, // sfix19_En18 
  input [18:0] Wgt_6_165, // sfix19_En18 
  input [18:0] Wgt_6_166, // sfix19_En18 
  input [18:0] Wgt_6_167, // sfix19_En18 
  input [18:0] Wgt_6_168, // sfix19_En18 
  input [18:0] Wgt_6_169, // sfix19_En18 
  input [18:0] Wgt_6_170, // sfix19_En18 
  input [18:0] Wgt_6_171, // sfix19_En18 
  input [18:0] Wgt_6_172, // sfix19_En18 
  input [18:0] Wgt_6_173, // sfix19_En18 
  input [18:0] Wgt_6_174, // sfix19_En18 
  input [18:0] Wgt_6_175, // sfix19_En18 
  input [18:0] Wgt_6_176, // sfix19_En18 
  input [18:0] Wgt_6_177, // sfix19_En18 
  input [18:0] Wgt_6_178, // sfix19_En18 
  input [18:0] Wgt_6_179, // sfix19_En18 
  input [18:0] Wgt_6_180, // sfix19_En18 
  input [18:0] Wgt_6_181, // sfix19_En18 
  input [18:0] Wgt_6_182, // sfix19_En18 
  input [18:0] Wgt_6_183, // sfix19_En18 
  input [18:0] Wgt_6_184, // sfix19_En18 
  input [18:0] Wgt_6_185, // sfix19_En18 
  input [18:0] Wgt_6_186, // sfix19_En18 
  input [18:0] Wgt_6_187, // sfix19_En18 
  input [18:0] Wgt_6_188, // sfix19_En18 
  input [18:0] Wgt_6_189, // sfix19_En18 
  input [18:0] Wgt_6_190, // sfix19_En18 
  input [18:0] Wgt_6_191, // sfix19_En18 
  input [18:0] Wgt_6_192, // sfix19_En18 
  input [18:0] Wgt_6_193, // sfix19_En18 
  input [18:0] Wgt_6_194, // sfix19_En18 
  input [18:0] Wgt_6_195, // sfix19_En18 
  input [18:0] Wgt_6_196, // sfix19_En18 
  input [18:0] Wgt_6_197, // sfix19_En18 
  input [18:0] Wgt_6_198, // sfix19_En18 
  input [18:0] Wgt_6_199, // sfix19_En18 
  input [18:0] Wgt_6_200, // sfix19_En18 
  input [18:0] Wgt_6_201, // sfix19_En18 
  input [18:0] Wgt_6_202, // sfix19_En18 
  input [18:0] Wgt_6_203, // sfix19_En18 
  input [18:0] Wgt_6_204, // sfix19_En18 
  input [18:0] Wgt_6_205, // sfix19_En18 
  input [18:0] Wgt_6_206, // sfix19_En18 
  input [18:0] Wgt_6_207, // sfix19_En18 
  input [18:0] Wgt_6_208, // sfix19_En18 
  input [18:0] Wgt_6_209, // sfix19_En18 
  input [18:0] Wgt_6_210, // sfix19_En18 
  input [18:0] Wgt_6_211, // sfix19_En18 
  input [18:0] Wgt_6_212, // sfix19_En18 
  input [18:0] Wgt_6_213, // sfix19_En18 
  input [18:0] Wgt_6_214, // sfix19_En18 
  input [18:0] Wgt_6_215, // sfix19_En18 
  input [18:0] Wgt_6_216, // sfix19_En18 
  input [18:0] Wgt_6_217, // sfix19_En18 
  input [18:0] Wgt_6_218, // sfix19_En18 
  input [18:0] Wgt_6_219, // sfix19_En18 
  input [18:0] Wgt_6_220, // sfix19_En18 
  input [18:0] Wgt_6_221, // sfix19_En18 
  input [18:0] Wgt_6_222, // sfix19_En18 
  input [18:0] Wgt_6_223, // sfix19_En18 
  input [18:0] Wgt_6_224, // sfix19_En18 
  input [18:0] Wgt_6_225, // sfix19_En18 
  input [18:0] Wgt_6_226, // sfix19_En18 
  input [18:0] Wgt_6_227, // sfix19_En18 
  input [18:0] Wgt_6_228, // sfix19_En18 
  input [18:0] Wgt_6_229, // sfix19_En18 
  input [18:0] Wgt_6_230, // sfix19_En18 
  input [18:0] Wgt_6_231, // sfix19_En18 
  input [18:0] Wgt_6_232, // sfix19_En18 
  input [18:0] Wgt_6_233, // sfix19_En18 
  input [18:0] Wgt_6_234, // sfix19_En18 
  input [18:0] Wgt_6_235, // sfix19_En18 
  input [18:0] Wgt_6_236, // sfix19_En18 
  input [18:0] Wgt_6_237, // sfix19_En18 
  input [18:0] Wgt_6_238, // sfix19_En18 
  input [18:0] Wgt_6_239, // sfix19_En18 
  input [18:0] Wgt_6_240, // sfix19_En18 
  input [18:0] Wgt_6_241, // sfix19_En18 
  input [18:0] Wgt_6_242, // sfix19_En18 
  input [18:0] Wgt_6_243, // sfix19_En18 
  input [18:0] Wgt_6_244, // sfix19_En18 
  input [18:0] Wgt_6_245, // sfix19_En18 
  input [18:0] Wgt_6_246, // sfix19_En18 
  input [18:0] Wgt_6_247, // sfix19_En18 
  input [18:0] Wgt_6_248, // sfix19_En18 
  input [18:0] Wgt_6_249, // sfix19_En18 
  input [18:0] Wgt_6_250, // sfix19_En18 
  input [18:0] Wgt_6_251, // sfix19_En18 
  input [18:0] Wgt_6_252, // sfix19_En18 
  input [18:0] Wgt_6_253, // sfix19_En18 
  input [18:0] Wgt_6_254, // sfix19_En18 
  input [18:0] Wgt_6_255, // sfix19_En18 
  input [18:0] Wgt_6_256, // sfix19_En18 
  input [18:0] Wgt_6_257, // sfix19_En18 
  input [18:0] Wgt_6_258, // sfix19_En18 
  input [18:0] Wgt_6_259, // sfix19_En18 
  input [18:0] Wgt_6_260, // sfix19_En18 
  input [18:0] Wgt_6_261, // sfix19_En18 
  input [18:0] Wgt_6_262, // sfix19_En18 
  input [18:0] Wgt_6_263, // sfix19_En18 
  input [18:0] Wgt_6_264, // sfix19_En18 
  input [18:0] Wgt_6_265, // sfix19_En18 
  input [18:0] Wgt_6_266, // sfix19_En18 
  input [18:0] Wgt_6_267, // sfix19_En18 
  input [18:0] Wgt_6_268, // sfix19_En18 
  input [18:0] Wgt_6_269, // sfix19_En18 
  input [18:0] Wgt_6_270, // sfix19_En18 
  input [18:0] Wgt_6_271, // sfix19_En18 
  input [18:0] Wgt_6_272, // sfix19_En18 
  input [18:0] Wgt_6_273, // sfix19_En18 
  input [18:0] Wgt_6_274, // sfix19_En18 
  input [18:0] Wgt_6_275, // sfix19_En18 
  input [18:0] Wgt_6_276, // sfix19_En18 
  input [18:0] Wgt_6_277, // sfix19_En18 
  input [18:0] Wgt_6_278, // sfix19_En18 
  input [18:0] Wgt_6_279, // sfix19_En18 
  input [18:0] Wgt_6_280, // sfix19_En18 
  input [18:0] Wgt_6_281, // sfix19_En18 
  input [18:0] Wgt_6_282, // sfix19_En18 
  input [18:0] Wgt_6_283, // sfix19_En18 
  input [18:0] Wgt_6_284, // sfix19_En18 
  input [18:0] Wgt_6_285, // sfix19_En18 
  input [18:0] Wgt_6_286, // sfix19_En18 
  input [18:0] Wgt_6_287, // sfix19_En18 
  input [18:0] Wgt_6_288, // sfix19_En18 
  input [18:0] Wgt_6_289, // sfix19_En18 
  input [18:0] Wgt_6_290, // sfix19_En18 
  input [18:0] Wgt_6_291, // sfix19_En18 
  input [18:0] Wgt_6_292, // sfix19_En18 
  input [18:0] Wgt_6_293, // sfix19_En18 
  input [18:0] Wgt_6_294, // sfix19_En18 
  input [18:0] Wgt_6_295, // sfix19_En18 
  input [18:0] Wgt_6_296, // sfix19_En18 
  input [18:0] Wgt_6_297, // sfix19_En18 
  input [18:0] Wgt_6_298, // sfix19_En18 
  input [18:0] Wgt_6_299, // sfix19_En18 
  input [18:0] Wgt_6_300, // sfix19_En18 
  input [18:0] Wgt_6_301, // sfix19_En18 
  input [18:0] Wgt_6_302, // sfix19_En18 
  input [18:0] Wgt_6_303, // sfix19_En18 
  input [18:0] Wgt_6_304, // sfix19_En18 
  input [18:0] Wgt_6_305, // sfix19_En18 
  input [18:0] Wgt_6_306, // sfix19_En18 
  input [18:0] Wgt_6_307, // sfix19_En18 
  input [18:0] Wgt_6_308, // sfix19_En18 
  input [18:0] Wgt_6_309, // sfix19_En18 
  input [18:0] Wgt_6_310, // sfix19_En18 
  input [18:0] Wgt_6_311, // sfix19_En18 
  input [18:0] Wgt_6_312, // sfix19_En18 
  input [18:0] Wgt_6_313, // sfix19_En18 
  input [18:0] Wgt_6_314, // sfix19_En18 
  input [18:0] Wgt_6_315, // sfix19_En18 
  input [18:0] Wgt_6_316, // sfix19_En18 
  input [18:0] Wgt_6_317, // sfix19_En18 
  input [18:0] Wgt_6_318, // sfix19_En18 
  input [18:0] Wgt_6_319, // sfix19_En18 
  input [18:0] Wgt_6_320, // sfix19_En18 
  input [18:0] Wgt_6_321, // sfix19_En18 
  input [18:0] Wgt_6_322, // sfix19_En18 
  input [18:0] Wgt_6_323, // sfix19_En18 
  input [18:0] Wgt_6_324, // sfix19_En18 
  input [18:0] Wgt_6_325, // sfix19_En18 
  input [18:0] Wgt_6_326, // sfix19_En18 
  input [18:0] Wgt_6_327, // sfix19_En18 
  input [18:0] Wgt_6_328, // sfix19_En18 
  input [18:0] Wgt_6_329, // sfix19_En18 
  input [18:0] Wgt_6_330, // sfix19_En18 
  input [18:0] Wgt_6_331, // sfix19_En18 
  input [18:0] Wgt_6_332, // sfix19_En18 
  input [18:0] Wgt_6_333, // sfix19_En18 
  input [18:0] Wgt_6_334, // sfix19_En18 
  input [18:0] Wgt_6_335, // sfix19_En18 
  input [18:0] Wgt_6_336, // sfix19_En18 
  input [18:0] Wgt_6_337, // sfix19_En18 
  input [18:0] Wgt_6_338, // sfix19_En18 
  input [18:0] Wgt_6_339, // sfix19_En18 
  input [18:0] Wgt_6_340, // sfix19_En18 
  input [18:0] Wgt_6_341, // sfix19_En18 
  input [18:0] Wgt_6_342, // sfix19_En18 
  input [18:0] Wgt_6_343, // sfix19_En18 
  input [18:0] Wgt_6_344, // sfix19_En18 
  input [18:0] Wgt_6_345, // sfix19_En18 
  input [18:0] Wgt_6_346, // sfix19_En18 
  input [18:0] Wgt_6_347, // sfix19_En18 
  input [18:0] Wgt_6_348, // sfix19_En18 
  input [18:0] Wgt_6_349, // sfix19_En18 
  input [18:0] Wgt_6_350, // sfix19_En18 
  input [18:0] Wgt_6_351, // sfix19_En18 
  input [18:0] Wgt_6_352, // sfix19_En18 
  input [18:0] Wgt_6_353, // sfix19_En18 
  input [18:0] Wgt_6_354, // sfix19_En18 
  input [18:0] Wgt_6_355, // sfix19_En18 
  input [18:0] Wgt_6_356, // sfix19_En18 
  input [18:0] Wgt_6_357, // sfix19_En18 
  input [18:0] Wgt_6_358, // sfix19_En18 
  input [18:0] Wgt_6_359, // sfix19_En18 
  input [18:0] Wgt_6_360, // sfix19_En18 
  input [18:0] Wgt_6_361, // sfix19_En18 
  input [18:0] Wgt_6_362, // sfix19_En18 
  input [18:0] Wgt_6_363, // sfix19_En18 
  input [18:0] Wgt_6_364, // sfix19_En18 
  input [18:0] Wgt_6_365, // sfix19_En18 
  input [18:0] Wgt_6_366, // sfix19_En18 
  input [18:0] Wgt_6_367, // sfix19_En18 
  input [18:0] Wgt_6_368, // sfix19_En18 
  input [18:0] Wgt_6_369, // sfix19_En18 
  input [18:0] Wgt_6_370, // sfix19_En18 
  input [18:0] Wgt_6_371, // sfix19_En18 
  input [18:0] Wgt_6_372, // sfix19_En18 
  input [18:0] Wgt_6_373, // sfix19_En18 
  input [18:0] Wgt_6_374, // sfix19_En18 
  input [18:0] Wgt_6_375, // sfix19_En18 
  input [18:0] Wgt_6_376, // sfix19_En18 
  input [18:0] Wgt_6_377, // sfix19_En18 
  input [18:0] Wgt_6_378, // sfix19_En18 
  input [18:0] Wgt_6_379, // sfix19_En18 
  input [18:0] Wgt_6_380, // sfix19_En18 
  input [18:0] Wgt_6_381, // sfix19_En18 
  input [18:0] Wgt_6_382, // sfix19_En18 
  input [18:0] Wgt_6_383, // sfix19_En18 
  input [18:0] Wgt_6_384, // sfix19_En18 
  input [18:0] Wgt_6_385, // sfix19_En18 
  input [18:0] Wgt_6_386, // sfix19_En18 
  input [18:0] Wgt_6_387, // sfix19_En18 
  input [18:0] Wgt_6_388, // sfix19_En18 
  input [18:0] Wgt_6_389, // sfix19_En18 
  input [18:0] Wgt_6_390, // sfix19_En18 
  input [18:0] Wgt_6_391, // sfix19_En18 
  input [18:0] Wgt_6_392, // sfix19_En18 
  input [18:0] Wgt_6_393, // sfix19_En18 
  input [18:0] Wgt_6_394, // sfix19_En18 
  input [18:0] Wgt_6_395, // sfix19_En18 
  input [18:0] Wgt_6_396, // sfix19_En18 
  input [18:0] Wgt_6_397, // sfix19_En18 
  input [18:0] Wgt_6_398, // sfix19_En18 
  input [18:0] Wgt_6_399, // sfix19_En18 
  input [18:0] Wgt_6_400, // sfix19_En18 
  input [18:0] Wgt_6_401, // sfix19_En18 
  input [18:0] Wgt_6_402, // sfix19_En18 
  input [18:0] Wgt_6_403, // sfix19_En18 
  input [18:0] Wgt_6_404, // sfix19_En18 
  input [18:0] Wgt_6_405, // sfix19_En18 
  input [18:0] Wgt_6_406, // sfix19_En18 
  input [18:0] Wgt_6_407, // sfix19_En18 
  input [18:0] Wgt_6_408, // sfix19_En18 
  input [18:0] Wgt_6_409, // sfix19_En18 
  input [18:0] Wgt_6_410, // sfix19_En18 
  input [18:0] Wgt_6_411, // sfix19_En18 
  input [18:0] Wgt_6_412, // sfix19_En18 
  input [18:0] Wgt_6_413, // sfix19_En18 
  input [18:0] Wgt_6_414, // sfix19_En18 
  input [18:0] Wgt_6_415, // sfix19_En18 
  input [18:0] Wgt_6_416, // sfix19_En18 
  input [18:0] Wgt_6_417, // sfix19_En18 
  input [18:0] Wgt_6_418, // sfix19_En18 
  input [18:0] Wgt_6_419, // sfix19_En18 
  input [18:0] Wgt_6_420, // sfix19_En18 
  input [18:0] Wgt_6_421, // sfix19_En18 
  input [18:0] Wgt_6_422, // sfix19_En18 
  input [18:0] Wgt_6_423, // sfix19_En18 
  input [18:0] Wgt_6_424, // sfix19_En18 
  input [18:0] Wgt_6_425, // sfix19_En18 
  input [18:0] Wgt_6_426, // sfix19_En18 
  input [18:0] Wgt_6_427, // sfix19_En18 
  input [18:0] Wgt_6_428, // sfix19_En18 
  input [18:0] Wgt_6_429, // sfix19_En18 
  input [18:0] Wgt_6_430, // sfix19_En18 
  input [18:0] Wgt_6_431, // sfix19_En18 
  input [18:0] Wgt_6_432, // sfix19_En18 
  input [18:0] Wgt_6_433, // sfix19_En18 
  input [18:0] Wgt_6_434, // sfix19_En18 
  input [18:0] Wgt_6_435, // sfix19_En18 
  input [18:0] Wgt_6_436, // sfix19_En18 
  input [18:0] Wgt_6_437, // sfix19_En18 
  input [18:0] Wgt_6_438, // sfix19_En18 
  input [18:0] Wgt_6_439, // sfix19_En18 
  input [18:0] Wgt_6_440, // sfix19_En18 
  input [18:0] Wgt_6_441, // sfix19_En18 
  input [18:0] Wgt_6_442, // sfix19_En18 
  input [18:0] Wgt_6_443, // sfix19_En18 
  input [18:0] Wgt_6_444, // sfix19_En18 
  input [18:0] Wgt_6_445, // sfix19_En18 
  input [18:0] Wgt_6_446, // sfix19_En18 
  input [18:0] Wgt_6_447, // sfix19_En18 
  input [18:0] Wgt_6_448, // sfix19_En18 
  input [18:0] Wgt_6_449, // sfix19_En18 
  input [18:0] Wgt_6_450, // sfix19_En18 
  input [18:0] Wgt_6_451, // sfix19_En18 
  input [18:0] Wgt_6_452, // sfix19_En18 
  input [18:0] Wgt_6_453, // sfix19_En18 
  input [18:0] Wgt_6_454, // sfix19_En18 
  input [18:0] Wgt_6_455, // sfix19_En18 
  input [18:0] Wgt_6_456, // sfix19_En18 
  input [18:0] Wgt_6_457, // sfix19_En18 
  input [18:0] Wgt_6_458, // sfix19_En18 
  input [18:0] Wgt_6_459, // sfix19_En18 
  input [18:0] Wgt_6_460, // sfix19_En18 
  input [18:0] Wgt_6_461, // sfix19_En18 
  input [18:0] Wgt_6_462, // sfix19_En18 
  input [18:0] Wgt_6_463, // sfix19_En18 
  input [18:0] Wgt_6_464, // sfix19_En18 
  input [18:0] Wgt_6_465, // sfix19_En18 
  input [18:0] Wgt_6_466, // sfix19_En18 
  input [18:0] Wgt_6_467, // sfix19_En18 
  input [18:0] Wgt_6_468, // sfix19_En18 
  input [18:0] Wgt_6_469, // sfix19_En18 
  input [18:0] Wgt_6_470, // sfix19_En18 
  input [18:0] Wgt_6_471, // sfix19_En18 
  input [18:0] Wgt_6_472, // sfix19_En18 
  input [18:0] Wgt_6_473, // sfix19_En18 
  input [18:0] Wgt_6_474, // sfix19_En18 
  input [18:0] Wgt_6_475, // sfix19_En18 
  input [18:0] Wgt_6_476, // sfix19_En18 
  input [18:0] Wgt_6_477, // sfix19_En18 
  input [18:0] Wgt_6_478, // sfix19_En18 
  input [18:0] Wgt_6_479, // sfix19_En18 
  input [18:0] Wgt_6_480, // sfix19_En18 
  input [18:0] Wgt_6_481, // sfix19_En18 
  input [18:0] Wgt_6_482, // sfix19_En18 
  input [18:0] Wgt_6_483, // sfix19_En18 
  input [18:0] Wgt_6_484, // sfix19_En18 
  input [18:0] Wgt_6_485, // sfix19_En18 
  input [18:0] Wgt_6_486, // sfix19_En18 
  input [18:0] Wgt_6_487, // sfix19_En18 
  input [18:0] Wgt_6_488, // sfix19_En18 
  input [18:0] Wgt_6_489, // sfix19_En18 
  input [18:0] Wgt_6_490, // sfix19_En18 
  input [18:0] Wgt_6_491, // sfix19_En18 
  input [18:0] Wgt_6_492, // sfix19_En18 
  input [18:0] Wgt_6_493, // sfix19_En18 
  input [18:0] Wgt_6_494, // sfix19_En18 
  input [18:0] Wgt_6_495, // sfix19_En18 
  input [18:0] Wgt_6_496, // sfix19_En18 
  input [18:0] Wgt_6_497, // sfix19_En18 
  input [18:0] Wgt_6_498, // sfix19_En18 
  input [18:0] Wgt_6_499, // sfix19_En18 
  input [18:0] Wgt_6_500, // sfix19_En18 
  input [18:0] Wgt_6_501, // sfix19_En18 
  input [18:0] Wgt_6_502, // sfix19_En18 
  input [18:0] Wgt_6_503, // sfix19_En18 
  input [18:0] Wgt_6_504, // sfix19_En18 
  input [18:0] Wgt_6_505, // sfix19_En18 
  input [18:0] Wgt_6_506, // sfix19_En18 
  input [18:0] Wgt_6_507, // sfix19_En18 
  input [18:0] Wgt_6_508, // sfix19_En18 
  input [18:0] Wgt_6_509, // sfix19_En18 
  input [18:0] Wgt_6_510, // sfix19_En18 
  input [18:0] Wgt_6_511, // sfix19_En18 
  input [18:0] Wgt_6_512, // sfix19_En18 
  input [18:0] Wgt_6_513, // sfix19_En18 
  input [18:0] Wgt_6_514, // sfix19_En18 
  input [18:0] Wgt_6_515, // sfix19_En18 
  input [18:0] Wgt_6_516, // sfix19_En18 
  input [18:0] Wgt_6_517, // sfix19_En18 
  input [18:0] Wgt_6_518, // sfix19_En18 
  input [18:0] Wgt_6_519, // sfix19_En18 
  input [18:0] Wgt_6_520, // sfix19_En18 
  input [18:0] Wgt_6_521, // sfix19_En18 
  input [18:0] Wgt_6_522, // sfix19_En18 
  input [18:0] Wgt_6_523, // sfix19_En18 
  input [18:0] Wgt_6_524, // sfix19_En18 
  input [18:0] Wgt_6_525, // sfix19_En18 
  input [18:0] Wgt_6_526, // sfix19_En18 
  input [18:0] Wgt_6_527, // sfix19_En18 
  input [18:0] Wgt_6_528, // sfix19_En18 
  input [18:0] Wgt_6_529, // sfix19_En18 
  input [18:0] Wgt_6_530, // sfix19_En18 
  input [18:0] Wgt_6_531, // sfix19_En18 
  input [18:0] Wgt_6_532, // sfix19_En18 
  input [18:0] Wgt_6_533, // sfix19_En18 
  input [18:0] Wgt_6_534, // sfix19_En18 
  input [18:0] Wgt_6_535, // sfix19_En18 
  input [18:0] Wgt_6_536, // sfix19_En18 
  input [18:0] Wgt_6_537, // sfix19_En18 
  input [18:0] Wgt_6_538, // sfix19_En18 
  input [18:0] Wgt_6_539, // sfix19_En18 
  input [18:0] Wgt_6_540, // sfix19_En18 
  input [18:0] Wgt_6_541, // sfix19_En18 
  input [18:0] Wgt_6_542, // sfix19_En18 
  input [18:0] Wgt_6_543, // sfix19_En18 
  input [18:0] Wgt_6_544, // sfix19_En18 
  input [18:0] Wgt_6_545, // sfix19_En18 
  input [18:0] Wgt_6_546, // sfix19_En18 
  input [18:0] Wgt_6_547, // sfix19_En18 
  input [18:0] Wgt_6_548, // sfix19_En18 
  input [18:0] Wgt_6_549, // sfix19_En18 
  input [18:0] Wgt_6_550, // sfix19_En18 
  input [18:0] Wgt_6_551, // sfix19_En18 
  input [18:0] Wgt_6_552, // sfix19_En18 
  input [18:0] Wgt_6_553, // sfix19_En18 
  input [18:0] Wgt_6_554, // sfix19_En18 
  input [18:0] Wgt_6_555, // sfix19_En18 
  input [18:0] Wgt_6_556, // sfix19_En18 
  input [18:0] Wgt_6_557, // sfix19_En18 
  input [18:0] Wgt_6_558, // sfix19_En18 
  input [18:0] Wgt_6_559, // sfix19_En18 
  input [18:0] Wgt_6_560, // sfix19_En18 
  input [18:0] Wgt_6_561, // sfix19_En18 
  input [18:0] Wgt_6_562, // sfix19_En18 
  input [18:0] Wgt_6_563, // sfix19_En18 
  input [18:0] Wgt_6_564, // sfix19_En18 
  input [18:0] Wgt_6_565, // sfix19_En18 
  input [18:0] Wgt_6_566, // sfix19_En18 
  input [18:0] Wgt_6_567, // sfix19_En18 
  input [18:0] Wgt_6_568, // sfix19_En18 
  input [18:0] Wgt_6_569, // sfix19_En18 
  input [18:0] Wgt_6_570, // sfix19_En18 
  input [18:0] Wgt_6_571, // sfix19_En18 
  input [18:0] Wgt_6_572, // sfix19_En18 
  input [18:0] Wgt_6_573, // sfix19_En18 
  input [18:0] Wgt_6_574, // sfix19_En18 
  input [18:0] Wgt_6_575, // sfix19_En18 
  input [18:0] Wgt_6_576, // sfix19_En18 
  input [18:0] Wgt_6_577, // sfix19_En18 
  input [18:0] Wgt_6_578, // sfix19_En18 
  input [18:0] Wgt_6_579, // sfix19_En18 
  input [18:0] Wgt_6_580, // sfix19_En18 
  input [18:0] Wgt_6_581, // sfix19_En18 
  input [18:0] Wgt_6_582, // sfix19_En18 
  input [18:0] Wgt_6_583, // sfix19_En18 
  input [18:0] Wgt_6_584, // sfix19_En18 
  input [18:0] Wgt_6_585, // sfix19_En18 
  input [18:0] Wgt_6_586, // sfix19_En18 
  input [18:0] Wgt_6_587, // sfix19_En18 
  input [18:0] Wgt_6_588, // sfix19_En18 
  input [18:0] Wgt_6_589, // sfix19_En18 
  input [18:0] Wgt_6_590, // sfix19_En18 
  input [18:0] Wgt_6_591, // sfix19_En18 
  input [18:0] Wgt_6_592, // sfix19_En18 
  input [18:0] Wgt_6_593, // sfix19_En18 
  input [18:0] Wgt_6_594, // sfix19_En18 
  input [18:0] Wgt_6_595, // sfix19_En18 
  input [18:0] Wgt_6_596, // sfix19_En18 
  input [18:0] Wgt_6_597, // sfix19_En18 
  input [18:0] Wgt_6_598, // sfix19_En18 
  input [18:0] Wgt_6_599, // sfix19_En18 
  input [18:0] Wgt_6_600, // sfix19_En18 
  input [18:0] Wgt_6_601, // sfix19_En18 
  input [18:0] Wgt_6_602, // sfix19_En18 
  input [18:0] Wgt_6_603, // sfix19_En18 
  input [18:0] Wgt_6_604, // sfix19_En18 
  input [18:0] Wgt_6_605, // sfix19_En18 
  input [18:0] Wgt_6_606, // sfix19_En18 
  input [18:0] Wgt_6_607, // sfix19_En18 
  input [18:0] Wgt_6_608, // sfix19_En18 
  input [18:0] Wgt_6_609, // sfix19_En18 
  input [18:0] Wgt_6_610, // sfix19_En18 
  input [18:0] Wgt_6_611, // sfix19_En18 
  input [18:0] Wgt_6_612, // sfix19_En18 
  input [18:0] Wgt_6_613, // sfix19_En18 
  input [18:0] Wgt_6_614, // sfix19_En18 
  input [18:0] Wgt_6_615, // sfix19_En18 
  input [18:0] Wgt_6_616, // sfix19_En18 
  input [18:0] Wgt_6_617, // sfix19_En18 
  input [18:0] Wgt_6_618, // sfix19_En18 
  input [18:0] Wgt_6_619, // sfix19_En18 
  input [18:0] Wgt_6_620, // sfix19_En18 
  input [18:0] Wgt_6_621, // sfix19_En18 
  input [18:0] Wgt_6_622, // sfix19_En18 
  input [18:0] Wgt_6_623, // sfix19_En18 
  input [18:0] Wgt_6_624, // sfix19_En18 
  input [18:0] Wgt_6_625, // sfix19_En18 
  input [18:0] Wgt_6_626, // sfix19_En18 
  input [18:0] Wgt_6_627, // sfix19_En18 
  input [18:0] Wgt_6_628, // sfix19_En18 
  input [18:0] Wgt_6_629, // sfix19_En18 
  input [18:0] Wgt_6_630, // sfix19_En18 
  input [18:0] Wgt_6_631, // sfix19_En18 
  input [18:0] Wgt_6_632, // sfix19_En18 
  input [18:0] Wgt_6_633, // sfix19_En18 
  input [18:0] Wgt_6_634, // sfix19_En18 
  input [18:0] Wgt_6_635, // sfix19_En18 
  input [18:0] Wgt_6_636, // sfix19_En18 
  input [18:0] Wgt_6_637, // sfix19_En18 
  input [18:0] Wgt_6_638, // sfix19_En18 
  input [18:0] Wgt_6_639, // sfix19_En18 
  input [18:0] Wgt_6_640, // sfix19_En18 
  input [18:0] Wgt_6_641, // sfix19_En18 
  input [18:0] Wgt_6_642, // sfix19_En18 
  input [18:0] Wgt_6_643, // sfix19_En18 
  input [18:0] Wgt_6_644, // sfix19_En18 
  input [18:0] Wgt_6_645, // sfix19_En18 
  input [18:0] Wgt_6_646, // sfix19_En18 
  input [18:0] Wgt_6_647, // sfix19_En18 
  input [18:0] Wgt_6_648, // sfix19_En18 
  input [18:0] Wgt_6_649, // sfix19_En18 
  input [18:0] Wgt_6_650, // sfix19_En18 
  input [18:0] Wgt_6_651, // sfix19_En18 
  input [18:0] Wgt_6_652, // sfix19_En18 
  input [18:0] Wgt_6_653, // sfix19_En18 
  input [18:0] Wgt_6_654, // sfix19_En18 
  input [18:0] Wgt_6_655, // sfix19_En18 
  input [18:0] Wgt_6_656, // sfix19_En18 
  input [18:0] Wgt_6_657, // sfix19_En18 
  input [18:0] Wgt_6_658, // sfix19_En18 
  input [18:0] Wgt_6_659, // sfix19_En18 
  input [18:0] Wgt_6_660, // sfix19_En18 
  input [18:0] Wgt_6_661, // sfix19_En18 
  input [18:0] Wgt_6_662, // sfix19_En18 
  input [18:0] Wgt_6_663, // sfix19_En18 
  input [18:0] Wgt_6_664, // sfix19_En18 
  input [18:0] Wgt_6_665, // sfix19_En18 
  input [18:0] Wgt_6_666, // sfix19_En18 
  input [18:0] Wgt_6_667, // sfix19_En18 
  input [18:0] Wgt_6_668, // sfix19_En18 
  input [18:0] Wgt_6_669, // sfix19_En18 
  input [18:0] Wgt_6_670, // sfix19_En18 
  input [18:0] Wgt_6_671, // sfix19_En18 
  input [18:0] Wgt_6_672, // sfix19_En18 
  input [18:0] Wgt_6_673, // sfix19_En18 
  input [18:0] Wgt_6_674, // sfix19_En18 
  input [18:0] Wgt_6_675, // sfix19_En18 
  input [18:0] Wgt_6_676, // sfix19_En18 
  input [18:0] Wgt_6_677, // sfix19_En18 
  input [18:0] Wgt_6_678, // sfix19_En18 
  input [18:0] Wgt_6_679, // sfix19_En18 
  input [18:0] Wgt_6_680, // sfix19_En18 
  input [18:0] Wgt_6_681, // sfix19_En18 
  input [18:0] Wgt_6_682, // sfix19_En18 
  input [18:0] Wgt_6_683, // sfix19_En18 
  input [18:0] Wgt_6_684, // sfix19_En18 
  input [18:0] Wgt_6_685, // sfix19_En18 
  input [18:0] Wgt_6_686, // sfix19_En18 
  input [18:0] Wgt_6_687, // sfix19_En18 
  input [18:0] Wgt_6_688, // sfix19_En18 
  input [18:0] Wgt_6_689, // sfix19_En18 
  input [18:0] Wgt_6_690, // sfix19_En18 
  input [18:0] Wgt_6_691, // sfix19_En18 
  input [18:0] Wgt_6_692, // sfix19_En18 
  input [18:0] Wgt_6_693, // sfix19_En18 
  input [18:0] Wgt_6_694, // sfix19_En18 
  input [18:0] Wgt_6_695, // sfix19_En18 
  input [18:0] Wgt_6_696, // sfix19_En18 
  input [18:0] Wgt_6_697, // sfix19_En18 
  input [18:0] Wgt_6_698, // sfix19_En18 
  input [18:0] Wgt_6_699, // sfix19_En18 
  input [18:0] Wgt_6_700, // sfix19_En18 
  input [18:0] Wgt_6_701, // sfix19_En18 
  input [18:0] Wgt_6_702, // sfix19_En18 
  input [18:0] Wgt_6_703, // sfix19_En18 
  input [18:0] Wgt_6_704, // sfix19_En18 
  input [18:0] Wgt_6_705, // sfix19_En18 
  input [18:0] Wgt_6_706, // sfix19_En18 
  input [18:0] Wgt_6_707, // sfix19_En18 
  input [18:0] Wgt_6_708, // sfix19_En18 
  input [18:0] Wgt_6_709, // sfix19_En18 
  input [18:0] Wgt_6_710, // sfix19_En18 
  input [18:0] Wgt_6_711, // sfix19_En18 
  input [18:0] Wgt_6_712, // sfix19_En18 
  input [18:0] Wgt_6_713, // sfix19_En18 
  input [18:0] Wgt_6_714, // sfix19_En18 
  input [18:0] Wgt_6_715, // sfix19_En18 
  input [18:0] Wgt_6_716, // sfix19_En18 
  input [18:0] Wgt_6_717, // sfix19_En18 
  input [18:0] Wgt_6_718, // sfix19_En18 
  input [18:0] Wgt_6_719, // sfix19_En18 
  input [18:0] Wgt_6_720, // sfix19_En18 
  input [18:0] Wgt_6_721, // sfix19_En18 
  input [18:0] Wgt_6_722, // sfix19_En18 
  input [18:0] Wgt_6_723, // sfix19_En18 
  input [18:0] Wgt_6_724, // sfix19_En18 
  input [18:0] Wgt_6_725, // sfix19_En18 
  input [18:0] Wgt_6_726, // sfix19_En18 
  input [18:0] Wgt_6_727, // sfix19_En18 
  input [18:0] Wgt_6_728, // sfix19_En18 
  input [18:0] Wgt_6_729, // sfix19_En18 
  input [18:0] Wgt_6_730, // sfix19_En18 
  input [18:0] Wgt_6_731, // sfix19_En18 
  input [18:0] Wgt_6_732, // sfix19_En18 
  input [18:0] Wgt_6_733, // sfix19_En18 
  input [18:0] Wgt_6_734, // sfix19_En18 
  input [18:0] Wgt_6_735, // sfix19_En18 
  input [18:0] Wgt_6_736, // sfix19_En18 
  input [18:0] Wgt_6_737, // sfix19_En18 
  input [18:0] Wgt_6_738, // sfix19_En18 
  input [18:0] Wgt_6_739, // sfix19_En18 
  input [18:0] Wgt_6_740, // sfix19_En18 
  input [18:0] Wgt_6_741, // sfix19_En18 
  input [18:0] Wgt_6_742, // sfix19_En18 
  input [18:0] Wgt_6_743, // sfix19_En18 
  input [18:0] Wgt_6_744, // sfix19_En18 
  input [18:0] Wgt_6_745, // sfix19_En18 
  input [18:0] Wgt_6_746, // sfix19_En18 
  input [18:0] Wgt_6_747, // sfix19_En18 
  input [18:0] Wgt_6_748, // sfix19_En18 
  input [18:0] Wgt_6_749, // sfix19_En18 
  input [18:0] Wgt_6_750, // sfix19_En18 
  input [18:0] Wgt_6_751, // sfix19_En18 
  input [18:0] Wgt_6_752, // sfix19_En18 
  input [18:0] Wgt_6_753, // sfix19_En18 
  input [18:0] Wgt_6_754, // sfix19_En18 
  input [18:0] Wgt_6_755, // sfix19_En18 
  input [18:0] Wgt_6_756, // sfix19_En18 
  input [18:0] Wgt_6_757, // sfix19_En18 
  input [18:0] Wgt_6_758, // sfix19_En18 
  input [18:0] Wgt_6_759, // sfix19_En18 
  input [18:0] Wgt_6_760, // sfix19_En18 
  input [18:0] Wgt_6_761, // sfix19_En18 
  input [18:0] Wgt_6_762, // sfix19_En18 
  input [18:0] Wgt_6_763, // sfix19_En18 
  input [18:0] Wgt_6_764, // sfix19_En18 
  input [18:0] Wgt_6_765, // sfix19_En18 
  input [18:0] Wgt_6_766, // sfix19_En18 
  input [18:0] Wgt_6_767, // sfix19_En18 
  input [18:0] Wgt_6_768, // sfix19_En18 
  input [18:0] Wgt_6_769, // sfix19_En18 
  input [18:0] Wgt_6_770, // sfix19_En18 
  input [18:0] Wgt_6_771, // sfix19_En18 
  input [18:0] Wgt_6_772, // sfix19_En18 
  input [18:0] Wgt_6_773, // sfix19_En18 
  input [18:0] Wgt_6_774, // sfix19_En18 
  input [18:0] Wgt_6_775, // sfix19_En18 
  input [18:0] Wgt_6_776, // sfix19_En18 
  input [18:0] Wgt_6_777, // sfix19_En18 
  input [18:0] Wgt_6_778, // sfix19_En18 
  input [18:0] Wgt_6_779, // sfix19_En18 
  input [18:0] Wgt_6_780, // sfix19_En18 
  input [18:0] Wgt_6_781, // sfix19_En18 
  input [18:0] Wgt_6_782, // sfix19_En18 
  input [18:0] Wgt_6_783, // sfix19_En18 
  input [18:0] Wgt_6_784, // sfix19_En18 
  input [18:0] Wgt_7_0, // sfix19_En18 
  input [18:0] Wgt_7_1, // sfix19_En18 
  input [18:0] Wgt_7_2, // sfix19_En18 
  input [18:0] Wgt_7_3, // sfix19_En18 
  input [18:0] Wgt_7_4, // sfix19_En18 
  input [18:0] Wgt_7_5, // sfix19_En18 
  input [18:0] Wgt_7_6, // sfix19_En18 
  input [18:0] Wgt_7_7, // sfix19_En18 
  input [18:0] Wgt_7_8, // sfix19_En18 
  input [18:0] Wgt_7_9, // sfix19_En18 
  input [18:0] Wgt_7_10, // sfix19_En18 
  input [18:0] Wgt_7_11, // sfix19_En18 
  input [18:0] Wgt_7_12, // sfix19_En18 
  input [18:0] Wgt_7_13, // sfix19_En18 
  input [18:0] Wgt_7_14, // sfix19_En18 
  input [18:0] Wgt_7_15, // sfix19_En18 
  input [18:0] Wgt_7_16, // sfix19_En18 
  input [18:0] Wgt_7_17, // sfix19_En18 
  input [18:0] Wgt_7_18, // sfix19_En18 
  input [18:0] Wgt_7_19, // sfix19_En18 
  input [18:0] Wgt_7_20, // sfix19_En18 
  input [18:0] Wgt_7_21, // sfix19_En18 
  input [18:0] Wgt_7_22, // sfix19_En18 
  input [18:0] Wgt_7_23, // sfix19_En18 
  input [18:0] Wgt_7_24, // sfix19_En18 
  input [18:0] Wgt_7_25, // sfix19_En18 
  input [18:0] Wgt_7_26, // sfix19_En18 
  input [18:0] Wgt_7_27, // sfix19_En18 
  input [18:0] Wgt_7_28, // sfix19_En18 
  input [18:0] Wgt_7_29, // sfix19_En18 
  input [18:0] Wgt_7_30, // sfix19_En18 
  input [18:0] Wgt_7_31, // sfix19_En18 
  input [18:0] Wgt_7_32, // sfix19_En18 
  input [18:0] Wgt_7_33, // sfix19_En18 
  input [18:0] Wgt_7_34, // sfix19_En18 
  input [18:0] Wgt_7_35, // sfix19_En18 
  input [18:0] Wgt_7_36, // sfix19_En18 
  input [18:0] Wgt_7_37, // sfix19_En18 
  input [18:0] Wgt_7_38, // sfix19_En18 
  input [18:0] Wgt_7_39, // sfix19_En18 
  input [18:0] Wgt_7_40, // sfix19_En18 
  input [18:0] Wgt_7_41, // sfix19_En18 
  input [18:0] Wgt_7_42, // sfix19_En18 
  input [18:0] Wgt_7_43, // sfix19_En18 
  input [18:0] Wgt_7_44, // sfix19_En18 
  input [18:0] Wgt_7_45, // sfix19_En18 
  input [18:0] Wgt_7_46, // sfix19_En18 
  input [18:0] Wgt_7_47, // sfix19_En18 
  input [18:0] Wgt_7_48, // sfix19_En18 
  input [18:0] Wgt_7_49, // sfix19_En18 
  input [18:0] Wgt_7_50, // sfix19_En18 
  input [18:0] Wgt_7_51, // sfix19_En18 
  input [18:0] Wgt_7_52, // sfix19_En18 
  input [18:0] Wgt_7_53, // sfix19_En18 
  input [18:0] Wgt_7_54, // sfix19_En18 
  input [18:0] Wgt_7_55, // sfix19_En18 
  input [18:0] Wgt_7_56, // sfix19_En18 
  input [18:0] Wgt_7_57, // sfix19_En18 
  input [18:0] Wgt_7_58, // sfix19_En18 
  input [18:0] Wgt_7_59, // sfix19_En18 
  input [18:0] Wgt_7_60, // sfix19_En18 
  input [18:0] Wgt_7_61, // sfix19_En18 
  input [18:0] Wgt_7_62, // sfix19_En18 
  input [18:0] Wgt_7_63, // sfix19_En18 
  input [18:0] Wgt_7_64, // sfix19_En18 
  input [18:0] Wgt_7_65, // sfix19_En18 
  input [18:0] Wgt_7_66, // sfix19_En18 
  input [18:0] Wgt_7_67, // sfix19_En18 
  input [18:0] Wgt_7_68, // sfix19_En18 
  input [18:0] Wgt_7_69, // sfix19_En18 
  input [18:0] Wgt_7_70, // sfix19_En18 
  input [18:0] Wgt_7_71, // sfix19_En18 
  input [18:0] Wgt_7_72, // sfix19_En18 
  input [18:0] Wgt_7_73, // sfix19_En18 
  input [18:0] Wgt_7_74, // sfix19_En18 
  input [18:0] Wgt_7_75, // sfix19_En18 
  input [18:0] Wgt_7_76, // sfix19_En18 
  input [18:0] Wgt_7_77, // sfix19_En18 
  input [18:0] Wgt_7_78, // sfix19_En18 
  input [18:0] Wgt_7_79, // sfix19_En18 
  input [18:0] Wgt_7_80, // sfix19_En18 
  input [18:0] Wgt_7_81, // sfix19_En18 
  input [18:0] Wgt_7_82, // sfix19_En18 
  input [18:0] Wgt_7_83, // sfix19_En18 
  input [18:0] Wgt_7_84, // sfix19_En18 
  input [18:0] Wgt_7_85, // sfix19_En18 
  input [18:0] Wgt_7_86, // sfix19_En18 
  input [18:0] Wgt_7_87, // sfix19_En18 
  input [18:0] Wgt_7_88, // sfix19_En18 
  input [18:0] Wgt_7_89, // sfix19_En18 
  input [18:0] Wgt_7_90, // sfix19_En18 
  input [18:0] Wgt_7_91, // sfix19_En18 
  input [18:0] Wgt_7_92, // sfix19_En18 
  input [18:0] Wgt_7_93, // sfix19_En18 
  input [18:0] Wgt_7_94, // sfix19_En18 
  input [18:0] Wgt_7_95, // sfix19_En18 
  input [18:0] Wgt_7_96, // sfix19_En18 
  input [18:0] Wgt_7_97, // sfix19_En18 
  input [18:0] Wgt_7_98, // sfix19_En18 
  input [18:0] Wgt_7_99, // sfix19_En18 
  input [18:0] Wgt_7_100, // sfix19_En18 
  input [18:0] Wgt_7_101, // sfix19_En18 
  input [18:0] Wgt_7_102, // sfix19_En18 
  input [18:0] Wgt_7_103, // sfix19_En18 
  input [18:0] Wgt_7_104, // sfix19_En18 
  input [18:0] Wgt_7_105, // sfix19_En18 
  input [18:0] Wgt_7_106, // sfix19_En18 
  input [18:0] Wgt_7_107, // sfix19_En18 
  input [18:0] Wgt_7_108, // sfix19_En18 
  input [18:0] Wgt_7_109, // sfix19_En18 
  input [18:0] Wgt_7_110, // sfix19_En18 
  input [18:0] Wgt_7_111, // sfix19_En18 
  input [18:0] Wgt_7_112, // sfix19_En18 
  input [18:0] Wgt_7_113, // sfix19_En18 
  input [18:0] Wgt_7_114, // sfix19_En18 
  input [18:0] Wgt_7_115, // sfix19_En18 
  input [18:0] Wgt_7_116, // sfix19_En18 
  input [18:0] Wgt_7_117, // sfix19_En18 
  input [18:0] Wgt_7_118, // sfix19_En18 
  input [18:0] Wgt_7_119, // sfix19_En18 
  input [18:0] Wgt_7_120, // sfix19_En18 
  input [18:0] Wgt_7_121, // sfix19_En18 
  input [18:0] Wgt_7_122, // sfix19_En18 
  input [18:0] Wgt_7_123, // sfix19_En18 
  input [18:0] Wgt_7_124, // sfix19_En18 
  input [18:0] Wgt_7_125, // sfix19_En18 
  input [18:0] Wgt_7_126, // sfix19_En18 
  input [18:0] Wgt_7_127, // sfix19_En18 
  input [18:0] Wgt_7_128, // sfix19_En18 
  input [18:0] Wgt_7_129, // sfix19_En18 
  input [18:0] Wgt_7_130, // sfix19_En18 
  input [18:0] Wgt_7_131, // sfix19_En18 
  input [18:0] Wgt_7_132, // sfix19_En18 
  input [18:0] Wgt_7_133, // sfix19_En18 
  input [18:0] Wgt_7_134, // sfix19_En18 
  input [18:0] Wgt_7_135, // sfix19_En18 
  input [18:0] Wgt_7_136, // sfix19_En18 
  input [18:0] Wgt_7_137, // sfix19_En18 
  input [18:0] Wgt_7_138, // sfix19_En18 
  input [18:0] Wgt_7_139, // sfix19_En18 
  input [18:0] Wgt_7_140, // sfix19_En18 
  input [18:0] Wgt_7_141, // sfix19_En18 
  input [18:0] Wgt_7_142, // sfix19_En18 
  input [18:0] Wgt_7_143, // sfix19_En18 
  input [18:0] Wgt_7_144, // sfix19_En18 
  input [18:0] Wgt_7_145, // sfix19_En18 
  input [18:0] Wgt_7_146, // sfix19_En18 
  input [18:0] Wgt_7_147, // sfix19_En18 
  input [18:0] Wgt_7_148, // sfix19_En18 
  input [18:0] Wgt_7_149, // sfix19_En18 
  input [18:0] Wgt_7_150, // sfix19_En18 
  input [18:0] Wgt_7_151, // sfix19_En18 
  input [18:0] Wgt_7_152, // sfix19_En18 
  input [18:0] Wgt_7_153, // sfix19_En18 
  input [18:0] Wgt_7_154, // sfix19_En18 
  input [18:0] Wgt_7_155, // sfix19_En18 
  input [18:0] Wgt_7_156, // sfix19_En18 
  input [18:0] Wgt_7_157, // sfix19_En18 
  input [18:0] Wgt_7_158, // sfix19_En18 
  input [18:0] Wgt_7_159, // sfix19_En18 
  input [18:0] Wgt_7_160, // sfix19_En18 
  input [18:0] Wgt_7_161, // sfix19_En18 
  input [18:0] Wgt_7_162, // sfix19_En18 
  input [18:0] Wgt_7_163, // sfix19_En18 
  input [18:0] Wgt_7_164, // sfix19_En18 
  input [18:0] Wgt_7_165, // sfix19_En18 
  input [18:0] Wgt_7_166, // sfix19_En18 
  input [18:0] Wgt_7_167, // sfix19_En18 
  input [18:0] Wgt_7_168, // sfix19_En18 
  input [18:0] Wgt_7_169, // sfix19_En18 
  input [18:0] Wgt_7_170, // sfix19_En18 
  input [18:0] Wgt_7_171, // sfix19_En18 
  input [18:0] Wgt_7_172, // sfix19_En18 
  input [18:0] Wgt_7_173, // sfix19_En18 
  input [18:0] Wgt_7_174, // sfix19_En18 
  input [18:0] Wgt_7_175, // sfix19_En18 
  input [18:0] Wgt_7_176, // sfix19_En18 
  input [18:0] Wgt_7_177, // sfix19_En18 
  input [18:0] Wgt_7_178, // sfix19_En18 
  input [18:0] Wgt_7_179, // sfix19_En18 
  input [18:0] Wgt_7_180, // sfix19_En18 
  input [18:0] Wgt_7_181, // sfix19_En18 
  input [18:0] Wgt_7_182, // sfix19_En18 
  input [18:0] Wgt_7_183, // sfix19_En18 
  input [18:0] Wgt_7_184, // sfix19_En18 
  input [18:0] Wgt_7_185, // sfix19_En18 
  input [18:0] Wgt_7_186, // sfix19_En18 
  input [18:0] Wgt_7_187, // sfix19_En18 
  input [18:0] Wgt_7_188, // sfix19_En18 
  input [18:0] Wgt_7_189, // sfix19_En18 
  input [18:0] Wgt_7_190, // sfix19_En18 
  input [18:0] Wgt_7_191, // sfix19_En18 
  input [18:0] Wgt_7_192, // sfix19_En18 
  input [18:0] Wgt_7_193, // sfix19_En18 
  input [18:0] Wgt_7_194, // sfix19_En18 
  input [18:0] Wgt_7_195, // sfix19_En18 
  input [18:0] Wgt_7_196, // sfix19_En18 
  input [18:0] Wgt_7_197, // sfix19_En18 
  input [18:0] Wgt_7_198, // sfix19_En18 
  input [18:0] Wgt_7_199, // sfix19_En18 
  input [18:0] Wgt_7_200, // sfix19_En18 
  input [18:0] Wgt_7_201, // sfix19_En18 
  input [18:0] Wgt_7_202, // sfix19_En18 
  input [18:0] Wgt_7_203, // sfix19_En18 
  input [18:0] Wgt_7_204, // sfix19_En18 
  input [18:0] Wgt_7_205, // sfix19_En18 
  input [18:0] Wgt_7_206, // sfix19_En18 
  input [18:0] Wgt_7_207, // sfix19_En18 
  input [18:0] Wgt_7_208, // sfix19_En18 
  input [18:0] Wgt_7_209, // sfix19_En18 
  input [18:0] Wgt_7_210, // sfix19_En18 
  input [18:0] Wgt_7_211, // sfix19_En18 
  input [18:0] Wgt_7_212, // sfix19_En18 
  input [18:0] Wgt_7_213, // sfix19_En18 
  input [18:0] Wgt_7_214, // sfix19_En18 
  input [18:0] Wgt_7_215, // sfix19_En18 
  input [18:0] Wgt_7_216, // sfix19_En18 
  input [18:0] Wgt_7_217, // sfix19_En18 
  input [18:0] Wgt_7_218, // sfix19_En18 
  input [18:0] Wgt_7_219, // sfix19_En18 
  input [18:0] Wgt_7_220, // sfix19_En18 
  input [18:0] Wgt_7_221, // sfix19_En18 
  input [18:0] Wgt_7_222, // sfix19_En18 
  input [18:0] Wgt_7_223, // sfix19_En18 
  input [18:0] Wgt_7_224, // sfix19_En18 
  input [18:0] Wgt_7_225, // sfix19_En18 
  input [18:0] Wgt_7_226, // sfix19_En18 
  input [18:0] Wgt_7_227, // sfix19_En18 
  input [18:0] Wgt_7_228, // sfix19_En18 
  input [18:0] Wgt_7_229, // sfix19_En18 
  input [18:0] Wgt_7_230, // sfix19_En18 
  input [18:0] Wgt_7_231, // sfix19_En18 
  input [18:0] Wgt_7_232, // sfix19_En18 
  input [18:0] Wgt_7_233, // sfix19_En18 
  input [18:0] Wgt_7_234, // sfix19_En18 
  input [18:0] Wgt_7_235, // sfix19_En18 
  input [18:0] Wgt_7_236, // sfix19_En18 
  input [18:0] Wgt_7_237, // sfix19_En18 
  input [18:0] Wgt_7_238, // sfix19_En18 
  input [18:0] Wgt_7_239, // sfix19_En18 
  input [18:0] Wgt_7_240, // sfix19_En18 
  input [18:0] Wgt_7_241, // sfix19_En18 
  input [18:0] Wgt_7_242, // sfix19_En18 
  input [18:0] Wgt_7_243, // sfix19_En18 
  input [18:0] Wgt_7_244, // sfix19_En18 
  input [18:0] Wgt_7_245, // sfix19_En18 
  input [18:0] Wgt_7_246, // sfix19_En18 
  input [18:0] Wgt_7_247, // sfix19_En18 
  input [18:0] Wgt_7_248, // sfix19_En18 
  input [18:0] Wgt_7_249, // sfix19_En18 
  input [18:0] Wgt_7_250, // sfix19_En18 
  input [18:0] Wgt_7_251, // sfix19_En18 
  input [18:0] Wgt_7_252, // sfix19_En18 
  input [18:0] Wgt_7_253, // sfix19_En18 
  input [18:0] Wgt_7_254, // sfix19_En18 
  input [18:0] Wgt_7_255, // sfix19_En18 
  input [18:0] Wgt_7_256, // sfix19_En18 
  input [18:0] Wgt_7_257, // sfix19_En18 
  input [18:0] Wgt_7_258, // sfix19_En18 
  input [18:0] Wgt_7_259, // sfix19_En18 
  input [18:0] Wgt_7_260, // sfix19_En18 
  input [18:0] Wgt_7_261, // sfix19_En18 
  input [18:0] Wgt_7_262, // sfix19_En18 
  input [18:0] Wgt_7_263, // sfix19_En18 
  input [18:0] Wgt_7_264, // sfix19_En18 
  input [18:0] Wgt_7_265, // sfix19_En18 
  input [18:0] Wgt_7_266, // sfix19_En18 
  input [18:0] Wgt_7_267, // sfix19_En18 
  input [18:0] Wgt_7_268, // sfix19_En18 
  input [18:0] Wgt_7_269, // sfix19_En18 
  input [18:0] Wgt_7_270, // sfix19_En18 
  input [18:0] Wgt_7_271, // sfix19_En18 
  input [18:0] Wgt_7_272, // sfix19_En18 
  input [18:0] Wgt_7_273, // sfix19_En18 
  input [18:0] Wgt_7_274, // sfix19_En18 
  input [18:0] Wgt_7_275, // sfix19_En18 
  input [18:0] Wgt_7_276, // sfix19_En18 
  input [18:0] Wgt_7_277, // sfix19_En18 
  input [18:0] Wgt_7_278, // sfix19_En18 
  input [18:0] Wgt_7_279, // sfix19_En18 
  input [18:0] Wgt_7_280, // sfix19_En18 
  input [18:0] Wgt_7_281, // sfix19_En18 
  input [18:0] Wgt_7_282, // sfix19_En18 
  input [18:0] Wgt_7_283, // sfix19_En18 
  input [18:0] Wgt_7_284, // sfix19_En18 
  input [18:0] Wgt_7_285, // sfix19_En18 
  input [18:0] Wgt_7_286, // sfix19_En18 
  input [18:0] Wgt_7_287, // sfix19_En18 
  input [18:0] Wgt_7_288, // sfix19_En18 
  input [18:0] Wgt_7_289, // sfix19_En18 
  input [18:0] Wgt_7_290, // sfix19_En18 
  input [18:0] Wgt_7_291, // sfix19_En18 
  input [18:0] Wgt_7_292, // sfix19_En18 
  input [18:0] Wgt_7_293, // sfix19_En18 
  input [18:0] Wgt_7_294, // sfix19_En18 
  input [18:0] Wgt_7_295, // sfix19_En18 
  input [18:0] Wgt_7_296, // sfix19_En18 
  input [18:0] Wgt_7_297, // sfix19_En18 
  input [18:0] Wgt_7_298, // sfix19_En18 
  input [18:0] Wgt_7_299, // sfix19_En18 
  input [18:0] Wgt_7_300, // sfix19_En18 
  input [18:0] Wgt_7_301, // sfix19_En18 
  input [18:0] Wgt_7_302, // sfix19_En18 
  input [18:0] Wgt_7_303, // sfix19_En18 
  input [18:0] Wgt_7_304, // sfix19_En18 
  input [18:0] Wgt_7_305, // sfix19_En18 
  input [18:0] Wgt_7_306, // sfix19_En18 
  input [18:0] Wgt_7_307, // sfix19_En18 
  input [18:0] Wgt_7_308, // sfix19_En18 
  input [18:0] Wgt_7_309, // sfix19_En18 
  input [18:0] Wgt_7_310, // sfix19_En18 
  input [18:0] Wgt_7_311, // sfix19_En18 
  input [18:0] Wgt_7_312, // sfix19_En18 
  input [18:0] Wgt_7_313, // sfix19_En18 
  input [18:0] Wgt_7_314, // sfix19_En18 
  input [18:0] Wgt_7_315, // sfix19_En18 
  input [18:0] Wgt_7_316, // sfix19_En18 
  input [18:0] Wgt_7_317, // sfix19_En18 
  input [18:0] Wgt_7_318, // sfix19_En18 
  input [18:0] Wgt_7_319, // sfix19_En18 
  input [18:0] Wgt_7_320, // sfix19_En18 
  input [18:0] Wgt_7_321, // sfix19_En18 
  input [18:0] Wgt_7_322, // sfix19_En18 
  input [18:0] Wgt_7_323, // sfix19_En18 
  input [18:0] Wgt_7_324, // sfix19_En18 
  input [18:0] Wgt_7_325, // sfix19_En18 
  input [18:0] Wgt_7_326, // sfix19_En18 
  input [18:0] Wgt_7_327, // sfix19_En18 
  input [18:0] Wgt_7_328, // sfix19_En18 
  input [18:0] Wgt_7_329, // sfix19_En18 
  input [18:0] Wgt_7_330, // sfix19_En18 
  input [18:0] Wgt_7_331, // sfix19_En18 
  input [18:0] Wgt_7_332, // sfix19_En18 
  input [18:0] Wgt_7_333, // sfix19_En18 
  input [18:0] Wgt_7_334, // sfix19_En18 
  input [18:0] Wgt_7_335, // sfix19_En18 
  input [18:0] Wgt_7_336, // sfix19_En18 
  input [18:0] Wgt_7_337, // sfix19_En18 
  input [18:0] Wgt_7_338, // sfix19_En18 
  input [18:0] Wgt_7_339, // sfix19_En18 
  input [18:0] Wgt_7_340, // sfix19_En18 
  input [18:0] Wgt_7_341, // sfix19_En18 
  input [18:0] Wgt_7_342, // sfix19_En18 
  input [18:0] Wgt_7_343, // sfix19_En18 
  input [18:0] Wgt_7_344, // sfix19_En18 
  input [18:0] Wgt_7_345, // sfix19_En18 
  input [18:0] Wgt_7_346, // sfix19_En18 
  input [18:0] Wgt_7_347, // sfix19_En18 
  input [18:0] Wgt_7_348, // sfix19_En18 
  input [18:0] Wgt_7_349, // sfix19_En18 
  input [18:0] Wgt_7_350, // sfix19_En18 
  input [18:0] Wgt_7_351, // sfix19_En18 
  input [18:0] Wgt_7_352, // sfix19_En18 
  input [18:0] Wgt_7_353, // sfix19_En18 
  input [18:0] Wgt_7_354, // sfix19_En18 
  input [18:0] Wgt_7_355, // sfix19_En18 
  input [18:0] Wgt_7_356, // sfix19_En18 
  input [18:0] Wgt_7_357, // sfix19_En18 
  input [18:0] Wgt_7_358, // sfix19_En18 
  input [18:0] Wgt_7_359, // sfix19_En18 
  input [18:0] Wgt_7_360, // sfix19_En18 
  input [18:0] Wgt_7_361, // sfix19_En18 
  input [18:0] Wgt_7_362, // sfix19_En18 
  input [18:0] Wgt_7_363, // sfix19_En18 
  input [18:0] Wgt_7_364, // sfix19_En18 
  input [18:0] Wgt_7_365, // sfix19_En18 
  input [18:0] Wgt_7_366, // sfix19_En18 
  input [18:0] Wgt_7_367, // sfix19_En18 
  input [18:0] Wgt_7_368, // sfix19_En18 
  input [18:0] Wgt_7_369, // sfix19_En18 
  input [18:0] Wgt_7_370, // sfix19_En18 
  input [18:0] Wgt_7_371, // sfix19_En18 
  input [18:0] Wgt_7_372, // sfix19_En18 
  input [18:0] Wgt_7_373, // sfix19_En18 
  input [18:0] Wgt_7_374, // sfix19_En18 
  input [18:0] Wgt_7_375, // sfix19_En18 
  input [18:0] Wgt_7_376, // sfix19_En18 
  input [18:0] Wgt_7_377, // sfix19_En18 
  input [18:0] Wgt_7_378, // sfix19_En18 
  input [18:0] Wgt_7_379, // sfix19_En18 
  input [18:0] Wgt_7_380, // sfix19_En18 
  input [18:0] Wgt_7_381, // sfix19_En18 
  input [18:0] Wgt_7_382, // sfix19_En18 
  input [18:0] Wgt_7_383, // sfix19_En18 
  input [18:0] Wgt_7_384, // sfix19_En18 
  input [18:0] Wgt_7_385, // sfix19_En18 
  input [18:0] Wgt_7_386, // sfix19_En18 
  input [18:0] Wgt_7_387, // sfix19_En18 
  input [18:0] Wgt_7_388, // sfix19_En18 
  input [18:0] Wgt_7_389, // sfix19_En18 
  input [18:0] Wgt_7_390, // sfix19_En18 
  input [18:0] Wgt_7_391, // sfix19_En18 
  input [18:0] Wgt_7_392, // sfix19_En18 
  input [18:0] Wgt_7_393, // sfix19_En18 
  input [18:0] Wgt_7_394, // sfix19_En18 
  input [18:0] Wgt_7_395, // sfix19_En18 
  input [18:0] Wgt_7_396, // sfix19_En18 
  input [18:0] Wgt_7_397, // sfix19_En18 
  input [18:0] Wgt_7_398, // sfix19_En18 
  input [18:0] Wgt_7_399, // sfix19_En18 
  input [18:0] Wgt_7_400, // sfix19_En18 
  input [18:0] Wgt_7_401, // sfix19_En18 
  input [18:0] Wgt_7_402, // sfix19_En18 
  input [18:0] Wgt_7_403, // sfix19_En18 
  input [18:0] Wgt_7_404, // sfix19_En18 
  input [18:0] Wgt_7_405, // sfix19_En18 
  input [18:0] Wgt_7_406, // sfix19_En18 
  input [18:0] Wgt_7_407, // sfix19_En18 
  input [18:0] Wgt_7_408, // sfix19_En18 
  input [18:0] Wgt_7_409, // sfix19_En18 
  input [18:0] Wgt_7_410, // sfix19_En18 
  input [18:0] Wgt_7_411, // sfix19_En18 
  input [18:0] Wgt_7_412, // sfix19_En18 
  input [18:0] Wgt_7_413, // sfix19_En18 
  input [18:0] Wgt_7_414, // sfix19_En18 
  input [18:0] Wgt_7_415, // sfix19_En18 
  input [18:0] Wgt_7_416, // sfix19_En18 
  input [18:0] Wgt_7_417, // sfix19_En18 
  input [18:0] Wgt_7_418, // sfix19_En18 
  input [18:0] Wgt_7_419, // sfix19_En18 
  input [18:0] Wgt_7_420, // sfix19_En18 
  input [18:0] Wgt_7_421, // sfix19_En18 
  input [18:0] Wgt_7_422, // sfix19_En18 
  input [18:0] Wgt_7_423, // sfix19_En18 
  input [18:0] Wgt_7_424, // sfix19_En18 
  input [18:0] Wgt_7_425, // sfix19_En18 
  input [18:0] Wgt_7_426, // sfix19_En18 
  input [18:0] Wgt_7_427, // sfix19_En18 
  input [18:0] Wgt_7_428, // sfix19_En18 
  input [18:0] Wgt_7_429, // sfix19_En18 
  input [18:0] Wgt_7_430, // sfix19_En18 
  input [18:0] Wgt_7_431, // sfix19_En18 
  input [18:0] Wgt_7_432, // sfix19_En18 
  input [18:0] Wgt_7_433, // sfix19_En18 
  input [18:0] Wgt_7_434, // sfix19_En18 
  input [18:0] Wgt_7_435, // sfix19_En18 
  input [18:0] Wgt_7_436, // sfix19_En18 
  input [18:0] Wgt_7_437, // sfix19_En18 
  input [18:0] Wgt_7_438, // sfix19_En18 
  input [18:0] Wgt_7_439, // sfix19_En18 
  input [18:0] Wgt_7_440, // sfix19_En18 
  input [18:0] Wgt_7_441, // sfix19_En18 
  input [18:0] Wgt_7_442, // sfix19_En18 
  input [18:0] Wgt_7_443, // sfix19_En18 
  input [18:0] Wgt_7_444, // sfix19_En18 
  input [18:0] Wgt_7_445, // sfix19_En18 
  input [18:0] Wgt_7_446, // sfix19_En18 
  input [18:0] Wgt_7_447, // sfix19_En18 
  input [18:0] Wgt_7_448, // sfix19_En18 
  input [18:0] Wgt_7_449, // sfix19_En18 
  input [18:0] Wgt_7_450, // sfix19_En18 
  input [18:0] Wgt_7_451, // sfix19_En18 
  input [18:0] Wgt_7_452, // sfix19_En18 
  input [18:0] Wgt_7_453, // sfix19_En18 
  input [18:0] Wgt_7_454, // sfix19_En18 
  input [18:0] Wgt_7_455, // sfix19_En18 
  input [18:0] Wgt_7_456, // sfix19_En18 
  input [18:0] Wgt_7_457, // sfix19_En18 
  input [18:0] Wgt_7_458, // sfix19_En18 
  input [18:0] Wgt_7_459, // sfix19_En18 
  input [18:0] Wgt_7_460, // sfix19_En18 
  input [18:0] Wgt_7_461, // sfix19_En18 
  input [18:0] Wgt_7_462, // sfix19_En18 
  input [18:0] Wgt_7_463, // sfix19_En18 
  input [18:0] Wgt_7_464, // sfix19_En18 
  input [18:0] Wgt_7_465, // sfix19_En18 
  input [18:0] Wgt_7_466, // sfix19_En18 
  input [18:0] Wgt_7_467, // sfix19_En18 
  input [18:0] Wgt_7_468, // sfix19_En18 
  input [18:0] Wgt_7_469, // sfix19_En18 
  input [18:0] Wgt_7_470, // sfix19_En18 
  input [18:0] Wgt_7_471, // sfix19_En18 
  input [18:0] Wgt_7_472, // sfix19_En18 
  input [18:0] Wgt_7_473, // sfix19_En18 
  input [18:0] Wgt_7_474, // sfix19_En18 
  input [18:0] Wgt_7_475, // sfix19_En18 
  input [18:0] Wgt_7_476, // sfix19_En18 
  input [18:0] Wgt_7_477, // sfix19_En18 
  input [18:0] Wgt_7_478, // sfix19_En18 
  input [18:0] Wgt_7_479, // sfix19_En18 
  input [18:0] Wgt_7_480, // sfix19_En18 
  input [18:0] Wgt_7_481, // sfix19_En18 
  input [18:0] Wgt_7_482, // sfix19_En18 
  input [18:0] Wgt_7_483, // sfix19_En18 
  input [18:0] Wgt_7_484, // sfix19_En18 
  input [18:0] Wgt_7_485, // sfix19_En18 
  input [18:0] Wgt_7_486, // sfix19_En18 
  input [18:0] Wgt_7_487, // sfix19_En18 
  input [18:0] Wgt_7_488, // sfix19_En18 
  input [18:0] Wgt_7_489, // sfix19_En18 
  input [18:0] Wgt_7_490, // sfix19_En18 
  input [18:0] Wgt_7_491, // sfix19_En18 
  input [18:0] Wgt_7_492, // sfix19_En18 
  input [18:0] Wgt_7_493, // sfix19_En18 
  input [18:0] Wgt_7_494, // sfix19_En18 
  input [18:0] Wgt_7_495, // sfix19_En18 
  input [18:0] Wgt_7_496, // sfix19_En18 
  input [18:0] Wgt_7_497, // sfix19_En18 
  input [18:0] Wgt_7_498, // sfix19_En18 
  input [18:0] Wgt_7_499, // sfix19_En18 
  input [18:0] Wgt_7_500, // sfix19_En18 
  input [18:0] Wgt_7_501, // sfix19_En18 
  input [18:0] Wgt_7_502, // sfix19_En18 
  input [18:0] Wgt_7_503, // sfix19_En18 
  input [18:0] Wgt_7_504, // sfix19_En18 
  input [18:0] Wgt_7_505, // sfix19_En18 
  input [18:0] Wgt_7_506, // sfix19_En18 
  input [18:0] Wgt_7_507, // sfix19_En18 
  input [18:0] Wgt_7_508, // sfix19_En18 
  input [18:0] Wgt_7_509, // sfix19_En18 
  input [18:0] Wgt_7_510, // sfix19_En18 
  input [18:0] Wgt_7_511, // sfix19_En18 
  input [18:0] Wgt_7_512, // sfix19_En18 
  input [18:0] Wgt_7_513, // sfix19_En18 
  input [18:0] Wgt_7_514, // sfix19_En18 
  input [18:0] Wgt_7_515, // sfix19_En18 
  input [18:0] Wgt_7_516, // sfix19_En18 
  input [18:0] Wgt_7_517, // sfix19_En18 
  input [18:0] Wgt_7_518, // sfix19_En18 
  input [18:0] Wgt_7_519, // sfix19_En18 
  input [18:0] Wgt_7_520, // sfix19_En18 
  input [18:0] Wgt_7_521, // sfix19_En18 
  input [18:0] Wgt_7_522, // sfix19_En18 
  input [18:0] Wgt_7_523, // sfix19_En18 
  input [18:0] Wgt_7_524, // sfix19_En18 
  input [18:0] Wgt_7_525, // sfix19_En18 
  input [18:0] Wgt_7_526, // sfix19_En18 
  input [18:0] Wgt_7_527, // sfix19_En18 
  input [18:0] Wgt_7_528, // sfix19_En18 
  input [18:0] Wgt_7_529, // sfix19_En18 
  input [18:0] Wgt_7_530, // sfix19_En18 
  input [18:0] Wgt_7_531, // sfix19_En18 
  input [18:0] Wgt_7_532, // sfix19_En18 
  input [18:0] Wgt_7_533, // sfix19_En18 
  input [18:0] Wgt_7_534, // sfix19_En18 
  input [18:0] Wgt_7_535, // sfix19_En18 
  input [18:0] Wgt_7_536, // sfix19_En18 
  input [18:0] Wgt_7_537, // sfix19_En18 
  input [18:0] Wgt_7_538, // sfix19_En18 
  input [18:0] Wgt_7_539, // sfix19_En18 
  input [18:0] Wgt_7_540, // sfix19_En18 
  input [18:0] Wgt_7_541, // sfix19_En18 
  input [18:0] Wgt_7_542, // sfix19_En18 
  input [18:0] Wgt_7_543, // sfix19_En18 
  input [18:0] Wgt_7_544, // sfix19_En18 
  input [18:0] Wgt_7_545, // sfix19_En18 
  input [18:0] Wgt_7_546, // sfix19_En18 
  input [18:0] Wgt_7_547, // sfix19_En18 
  input [18:0] Wgt_7_548, // sfix19_En18 
  input [18:0] Wgt_7_549, // sfix19_En18 
  input [18:0] Wgt_7_550, // sfix19_En18 
  input [18:0] Wgt_7_551, // sfix19_En18 
  input [18:0] Wgt_7_552, // sfix19_En18 
  input [18:0] Wgt_7_553, // sfix19_En18 
  input [18:0] Wgt_7_554, // sfix19_En18 
  input [18:0] Wgt_7_555, // sfix19_En18 
  input [18:0] Wgt_7_556, // sfix19_En18 
  input [18:0] Wgt_7_557, // sfix19_En18 
  input [18:0] Wgt_7_558, // sfix19_En18 
  input [18:0] Wgt_7_559, // sfix19_En18 
  input [18:0] Wgt_7_560, // sfix19_En18 
  input [18:0] Wgt_7_561, // sfix19_En18 
  input [18:0] Wgt_7_562, // sfix19_En18 
  input [18:0] Wgt_7_563, // sfix19_En18 
  input [18:0] Wgt_7_564, // sfix19_En18 
  input [18:0] Wgt_7_565, // sfix19_En18 
  input [18:0] Wgt_7_566, // sfix19_En18 
  input [18:0] Wgt_7_567, // sfix19_En18 
  input [18:0] Wgt_7_568, // sfix19_En18 
  input [18:0] Wgt_7_569, // sfix19_En18 
  input [18:0] Wgt_7_570, // sfix19_En18 
  input [18:0] Wgt_7_571, // sfix19_En18 
  input [18:0] Wgt_7_572, // sfix19_En18 
  input [18:0] Wgt_7_573, // sfix19_En18 
  input [18:0] Wgt_7_574, // sfix19_En18 
  input [18:0] Wgt_7_575, // sfix19_En18 
  input [18:0] Wgt_7_576, // sfix19_En18 
  input [18:0] Wgt_7_577, // sfix19_En18 
  input [18:0] Wgt_7_578, // sfix19_En18 
  input [18:0] Wgt_7_579, // sfix19_En18 
  input [18:0] Wgt_7_580, // sfix19_En18 
  input [18:0] Wgt_7_581, // sfix19_En18 
  input [18:0] Wgt_7_582, // sfix19_En18 
  input [18:0] Wgt_7_583, // sfix19_En18 
  input [18:0] Wgt_7_584, // sfix19_En18 
  input [18:0] Wgt_7_585, // sfix19_En18 
  input [18:0] Wgt_7_586, // sfix19_En18 
  input [18:0] Wgt_7_587, // sfix19_En18 
  input [18:0] Wgt_7_588, // sfix19_En18 
  input [18:0] Wgt_7_589, // sfix19_En18 
  input [18:0] Wgt_7_590, // sfix19_En18 
  input [18:0] Wgt_7_591, // sfix19_En18 
  input [18:0] Wgt_7_592, // sfix19_En18 
  input [18:0] Wgt_7_593, // sfix19_En18 
  input [18:0] Wgt_7_594, // sfix19_En18 
  input [18:0] Wgt_7_595, // sfix19_En18 
  input [18:0] Wgt_7_596, // sfix19_En18 
  input [18:0] Wgt_7_597, // sfix19_En18 
  input [18:0] Wgt_7_598, // sfix19_En18 
  input [18:0] Wgt_7_599, // sfix19_En18 
  input [18:0] Wgt_7_600, // sfix19_En18 
  input [18:0] Wgt_7_601, // sfix19_En18 
  input [18:0] Wgt_7_602, // sfix19_En18 
  input [18:0] Wgt_7_603, // sfix19_En18 
  input [18:0] Wgt_7_604, // sfix19_En18 
  input [18:0] Wgt_7_605, // sfix19_En18 
  input [18:0] Wgt_7_606, // sfix19_En18 
  input [18:0] Wgt_7_607, // sfix19_En18 
  input [18:0] Wgt_7_608, // sfix19_En18 
  input [18:0] Wgt_7_609, // sfix19_En18 
  input [18:0] Wgt_7_610, // sfix19_En18 
  input [18:0] Wgt_7_611, // sfix19_En18 
  input [18:0] Wgt_7_612, // sfix19_En18 
  input [18:0] Wgt_7_613, // sfix19_En18 
  input [18:0] Wgt_7_614, // sfix19_En18 
  input [18:0] Wgt_7_615, // sfix19_En18 
  input [18:0] Wgt_7_616, // sfix19_En18 
  input [18:0] Wgt_7_617, // sfix19_En18 
  input [18:0] Wgt_7_618, // sfix19_En18 
  input [18:0] Wgt_7_619, // sfix19_En18 
  input [18:0] Wgt_7_620, // sfix19_En18 
  input [18:0] Wgt_7_621, // sfix19_En18 
  input [18:0] Wgt_7_622, // sfix19_En18 
  input [18:0] Wgt_7_623, // sfix19_En18 
  input [18:0] Wgt_7_624, // sfix19_En18 
  input [18:0] Wgt_7_625, // sfix19_En18 
  input [18:0] Wgt_7_626, // sfix19_En18 
  input [18:0] Wgt_7_627, // sfix19_En18 
  input [18:0] Wgt_7_628, // sfix19_En18 
  input [18:0] Wgt_7_629, // sfix19_En18 
  input [18:0] Wgt_7_630, // sfix19_En18 
  input [18:0] Wgt_7_631, // sfix19_En18 
  input [18:0] Wgt_7_632, // sfix19_En18 
  input [18:0] Wgt_7_633, // sfix19_En18 
  input [18:0] Wgt_7_634, // sfix19_En18 
  input [18:0] Wgt_7_635, // sfix19_En18 
  input [18:0] Wgt_7_636, // sfix19_En18 
  input [18:0] Wgt_7_637, // sfix19_En18 
  input [18:0] Wgt_7_638, // sfix19_En18 
  input [18:0] Wgt_7_639, // sfix19_En18 
  input [18:0] Wgt_7_640, // sfix19_En18 
  input [18:0] Wgt_7_641, // sfix19_En18 
  input [18:0] Wgt_7_642, // sfix19_En18 
  input [18:0] Wgt_7_643, // sfix19_En18 
  input [18:0] Wgt_7_644, // sfix19_En18 
  input [18:0] Wgt_7_645, // sfix19_En18 
  input [18:0] Wgt_7_646, // sfix19_En18 
  input [18:0] Wgt_7_647, // sfix19_En18 
  input [18:0] Wgt_7_648, // sfix19_En18 
  input [18:0] Wgt_7_649, // sfix19_En18 
  input [18:0] Wgt_7_650, // sfix19_En18 
  input [18:0] Wgt_7_651, // sfix19_En18 
  input [18:0] Wgt_7_652, // sfix19_En18 
  input [18:0] Wgt_7_653, // sfix19_En18 
  input [18:0] Wgt_7_654, // sfix19_En18 
  input [18:0] Wgt_7_655, // sfix19_En18 
  input [18:0] Wgt_7_656, // sfix19_En18 
  input [18:0] Wgt_7_657, // sfix19_En18 
  input [18:0] Wgt_7_658, // sfix19_En18 
  input [18:0] Wgt_7_659, // sfix19_En18 
  input [18:0] Wgt_7_660, // sfix19_En18 
  input [18:0] Wgt_7_661, // sfix19_En18 
  input [18:0] Wgt_7_662, // sfix19_En18 
  input [18:0] Wgt_7_663, // sfix19_En18 
  input [18:0] Wgt_7_664, // sfix19_En18 
  input [18:0] Wgt_7_665, // sfix19_En18 
  input [18:0] Wgt_7_666, // sfix19_En18 
  input [18:0] Wgt_7_667, // sfix19_En18 
  input [18:0] Wgt_7_668, // sfix19_En18 
  input [18:0] Wgt_7_669, // sfix19_En18 
  input [18:0] Wgt_7_670, // sfix19_En18 
  input [18:0] Wgt_7_671, // sfix19_En18 
  input [18:0] Wgt_7_672, // sfix19_En18 
  input [18:0] Wgt_7_673, // sfix19_En18 
  input [18:0] Wgt_7_674, // sfix19_En18 
  input [18:0] Wgt_7_675, // sfix19_En18 
  input [18:0] Wgt_7_676, // sfix19_En18 
  input [18:0] Wgt_7_677, // sfix19_En18 
  input [18:0] Wgt_7_678, // sfix19_En18 
  input [18:0] Wgt_7_679, // sfix19_En18 
  input [18:0] Wgt_7_680, // sfix19_En18 
  input [18:0] Wgt_7_681, // sfix19_En18 
  input [18:0] Wgt_7_682, // sfix19_En18 
  input [18:0] Wgt_7_683, // sfix19_En18 
  input [18:0] Wgt_7_684, // sfix19_En18 
  input [18:0] Wgt_7_685, // sfix19_En18 
  input [18:0] Wgt_7_686, // sfix19_En18 
  input [18:0] Wgt_7_687, // sfix19_En18 
  input [18:0] Wgt_7_688, // sfix19_En18 
  input [18:0] Wgt_7_689, // sfix19_En18 
  input [18:0] Wgt_7_690, // sfix19_En18 
  input [18:0] Wgt_7_691, // sfix19_En18 
  input [18:0] Wgt_7_692, // sfix19_En18 
  input [18:0] Wgt_7_693, // sfix19_En18 
  input [18:0] Wgt_7_694, // sfix19_En18 
  input [18:0] Wgt_7_695, // sfix19_En18 
  input [18:0] Wgt_7_696, // sfix19_En18 
  input [18:0] Wgt_7_697, // sfix19_En18 
  input [18:0] Wgt_7_698, // sfix19_En18 
  input [18:0] Wgt_7_699, // sfix19_En18 
  input [18:0] Wgt_7_700, // sfix19_En18 
  input [18:0] Wgt_7_701, // sfix19_En18 
  input [18:0] Wgt_7_702, // sfix19_En18 
  input [18:0] Wgt_7_703, // sfix19_En18 
  input [18:0] Wgt_7_704, // sfix19_En18 
  input [18:0] Wgt_7_705, // sfix19_En18 
  input [18:0] Wgt_7_706, // sfix19_En18 
  input [18:0] Wgt_7_707, // sfix19_En18 
  input [18:0] Wgt_7_708, // sfix19_En18 
  input [18:0] Wgt_7_709, // sfix19_En18 
  input [18:0] Wgt_7_710, // sfix19_En18 
  input [18:0] Wgt_7_711, // sfix19_En18 
  input [18:0] Wgt_7_712, // sfix19_En18 
  input [18:0] Wgt_7_713, // sfix19_En18 
  input [18:0] Wgt_7_714, // sfix19_En18 
  input [18:0] Wgt_7_715, // sfix19_En18 
  input [18:0] Wgt_7_716, // sfix19_En18 
  input [18:0] Wgt_7_717, // sfix19_En18 
  input [18:0] Wgt_7_718, // sfix19_En18 
  input [18:0] Wgt_7_719, // sfix19_En18 
  input [18:0] Wgt_7_720, // sfix19_En18 
  input [18:0] Wgt_7_721, // sfix19_En18 
  input [18:0] Wgt_7_722, // sfix19_En18 
  input [18:0] Wgt_7_723, // sfix19_En18 
  input [18:0] Wgt_7_724, // sfix19_En18 
  input [18:0] Wgt_7_725, // sfix19_En18 
  input [18:0] Wgt_7_726, // sfix19_En18 
  input [18:0] Wgt_7_727, // sfix19_En18 
  input [18:0] Wgt_7_728, // sfix19_En18 
  input [18:0] Wgt_7_729, // sfix19_En18 
  input [18:0] Wgt_7_730, // sfix19_En18 
  input [18:0] Wgt_7_731, // sfix19_En18 
  input [18:0] Wgt_7_732, // sfix19_En18 
  input [18:0] Wgt_7_733, // sfix19_En18 
  input [18:0] Wgt_7_734, // sfix19_En18 
  input [18:0] Wgt_7_735, // sfix19_En18 
  input [18:0] Wgt_7_736, // sfix19_En18 
  input [18:0] Wgt_7_737, // sfix19_En18 
  input [18:0] Wgt_7_738, // sfix19_En18 
  input [18:0] Wgt_7_739, // sfix19_En18 
  input [18:0] Wgt_7_740, // sfix19_En18 
  input [18:0] Wgt_7_741, // sfix19_En18 
  input [18:0] Wgt_7_742, // sfix19_En18 
  input [18:0] Wgt_7_743, // sfix19_En18 
  input [18:0] Wgt_7_744, // sfix19_En18 
  input [18:0] Wgt_7_745, // sfix19_En18 
  input [18:0] Wgt_7_746, // sfix19_En18 
  input [18:0] Wgt_7_747, // sfix19_En18 
  input [18:0] Wgt_7_748, // sfix19_En18 
  input [18:0] Wgt_7_749, // sfix19_En18 
  input [18:0] Wgt_7_750, // sfix19_En18 
  input [18:0] Wgt_7_751, // sfix19_En18 
  input [18:0] Wgt_7_752, // sfix19_En18 
  input [18:0] Wgt_7_753, // sfix19_En18 
  input [18:0] Wgt_7_754, // sfix19_En18 
  input [18:0] Wgt_7_755, // sfix19_En18 
  input [18:0] Wgt_7_756, // sfix19_En18 
  input [18:0] Wgt_7_757, // sfix19_En18 
  input [18:0] Wgt_7_758, // sfix19_En18 
  input [18:0] Wgt_7_759, // sfix19_En18 
  input [18:0] Wgt_7_760, // sfix19_En18 
  input [18:0] Wgt_7_761, // sfix19_En18 
  input [18:0] Wgt_7_762, // sfix19_En18 
  input [18:0] Wgt_7_763, // sfix19_En18 
  input [18:0] Wgt_7_764, // sfix19_En18 
  input [18:0] Wgt_7_765, // sfix19_En18 
  input [18:0] Wgt_7_766, // sfix19_En18 
  input [18:0] Wgt_7_767, // sfix19_En18 
  input [18:0] Wgt_7_768, // sfix19_En18 
  input [18:0] Wgt_7_769, // sfix19_En18 
  input [18:0] Wgt_7_770, // sfix19_En18 
  input [18:0] Wgt_7_771, // sfix19_En18 
  input [18:0] Wgt_7_772, // sfix19_En18 
  input [18:0] Wgt_7_773, // sfix19_En18 
  input [18:0] Wgt_7_774, // sfix19_En18 
  input [18:0] Wgt_7_775, // sfix19_En18 
  input [18:0] Wgt_7_776, // sfix19_En18 
  input [18:0] Wgt_7_777, // sfix19_En18 
  input [18:0] Wgt_7_778, // sfix19_En18 
  input [18:0] Wgt_7_779, // sfix19_En18 
  input [18:0] Wgt_7_780, // sfix19_En18 
  input [18:0] Wgt_7_781, // sfix19_En18 
  input [18:0] Wgt_7_782, // sfix19_En18 
  input [18:0] Wgt_7_783, // sfix19_En18 
  input [18:0] Wgt_7_784, // sfix19_En18 
  input [18:0] Wgt_8_0, // sfix19_En18 
  input [18:0] Wgt_8_1, // sfix19_En18 
  input [18:0] Wgt_8_2, // sfix19_En18 
  input [18:0] Wgt_8_3, // sfix19_En18 
  input [18:0] Wgt_8_4, // sfix19_En18 
  input [18:0] Wgt_8_5, // sfix19_En18 
  input [18:0] Wgt_8_6, // sfix19_En18 
  input [18:0] Wgt_8_7, // sfix19_En18 
  input [18:0] Wgt_8_8, // sfix19_En18 
  input [18:0] Wgt_8_9, // sfix19_En18 
  input [18:0] Wgt_8_10, // sfix19_En18 
  input [18:0] Wgt_8_11, // sfix19_En18 
  input [18:0] Wgt_8_12, // sfix19_En18 
  input [18:0] Wgt_8_13, // sfix19_En18 
  input [18:0] Wgt_8_14, // sfix19_En18 
  input [18:0] Wgt_8_15, // sfix19_En18 
  input [18:0] Wgt_8_16, // sfix19_En18 
  input [18:0] Wgt_8_17, // sfix19_En18 
  input [18:0] Wgt_8_18, // sfix19_En18 
  input [18:0] Wgt_8_19, // sfix19_En18 
  input [18:0] Wgt_8_20, // sfix19_En18 
  input [18:0] Wgt_8_21, // sfix19_En18 
  input [18:0] Wgt_8_22, // sfix19_En18 
  input [18:0] Wgt_8_23, // sfix19_En18 
  input [18:0] Wgt_8_24, // sfix19_En18 
  input [18:0] Wgt_8_25, // sfix19_En18 
  input [18:0] Wgt_8_26, // sfix19_En18 
  input [18:0] Wgt_8_27, // sfix19_En18 
  input [18:0] Wgt_8_28, // sfix19_En18 
  input [18:0] Wgt_8_29, // sfix19_En18 
  input [18:0] Wgt_8_30, // sfix19_En18 
  input [18:0] Wgt_8_31, // sfix19_En18 
  input [18:0] Wgt_8_32, // sfix19_En18 
  input [18:0] Wgt_8_33, // sfix19_En18 
  input [18:0] Wgt_8_34, // sfix19_En18 
  input [18:0] Wgt_8_35, // sfix19_En18 
  input [18:0] Wgt_8_36, // sfix19_En18 
  input [18:0] Wgt_8_37, // sfix19_En18 
  input [18:0] Wgt_8_38, // sfix19_En18 
  input [18:0] Wgt_8_39, // sfix19_En18 
  input [18:0] Wgt_8_40, // sfix19_En18 
  input [18:0] Wgt_8_41, // sfix19_En18 
  input [18:0] Wgt_8_42, // sfix19_En18 
  input [18:0] Wgt_8_43, // sfix19_En18 
  input [18:0] Wgt_8_44, // sfix19_En18 
  input [18:0] Wgt_8_45, // sfix19_En18 
  input [18:0] Wgt_8_46, // sfix19_En18 
  input [18:0] Wgt_8_47, // sfix19_En18 
  input [18:0] Wgt_8_48, // sfix19_En18 
  input [18:0] Wgt_8_49, // sfix19_En18 
  input [18:0] Wgt_8_50, // sfix19_En18 
  input [18:0] Wgt_8_51, // sfix19_En18 
  input [18:0] Wgt_8_52, // sfix19_En18 
  input [18:0] Wgt_8_53, // sfix19_En18 
  input [18:0] Wgt_8_54, // sfix19_En18 
  input [18:0] Wgt_8_55, // sfix19_En18 
  input [18:0] Wgt_8_56, // sfix19_En18 
  input [18:0] Wgt_8_57, // sfix19_En18 
  input [18:0] Wgt_8_58, // sfix19_En18 
  input [18:0] Wgt_8_59, // sfix19_En18 
  input [18:0] Wgt_8_60, // sfix19_En18 
  input [18:0] Wgt_8_61, // sfix19_En18 
  input [18:0] Wgt_8_62, // sfix19_En18 
  input [18:0] Wgt_8_63, // sfix19_En18 
  input [18:0] Wgt_8_64, // sfix19_En18 
  input [18:0] Wgt_8_65, // sfix19_En18 
  input [18:0] Wgt_8_66, // sfix19_En18 
  input [18:0] Wgt_8_67, // sfix19_En18 
  input [18:0] Wgt_8_68, // sfix19_En18 
  input [18:0] Wgt_8_69, // sfix19_En18 
  input [18:0] Wgt_8_70, // sfix19_En18 
  input [18:0] Wgt_8_71, // sfix19_En18 
  input [18:0] Wgt_8_72, // sfix19_En18 
  input [18:0] Wgt_8_73, // sfix19_En18 
  input [18:0] Wgt_8_74, // sfix19_En18 
  input [18:0] Wgt_8_75, // sfix19_En18 
  input [18:0] Wgt_8_76, // sfix19_En18 
  input [18:0] Wgt_8_77, // sfix19_En18 
  input [18:0] Wgt_8_78, // sfix19_En18 
  input [18:0] Wgt_8_79, // sfix19_En18 
  input [18:0] Wgt_8_80, // sfix19_En18 
  input [18:0] Wgt_8_81, // sfix19_En18 
  input [18:0] Wgt_8_82, // sfix19_En18 
  input [18:0] Wgt_8_83, // sfix19_En18 
  input [18:0] Wgt_8_84, // sfix19_En18 
  input [18:0] Wgt_8_85, // sfix19_En18 
  input [18:0] Wgt_8_86, // sfix19_En18 
  input [18:0] Wgt_8_87, // sfix19_En18 
  input [18:0] Wgt_8_88, // sfix19_En18 
  input [18:0] Wgt_8_89, // sfix19_En18 
  input [18:0] Wgt_8_90, // sfix19_En18 
  input [18:0] Wgt_8_91, // sfix19_En18 
  input [18:0] Wgt_8_92, // sfix19_En18 
  input [18:0] Wgt_8_93, // sfix19_En18 
  input [18:0] Wgt_8_94, // sfix19_En18 
  input [18:0] Wgt_8_95, // sfix19_En18 
  input [18:0] Wgt_8_96, // sfix19_En18 
  input [18:0] Wgt_8_97, // sfix19_En18 
  input [18:0] Wgt_8_98, // sfix19_En18 
  input [18:0] Wgt_8_99, // sfix19_En18 
  input [18:0] Wgt_8_100, // sfix19_En18 
  input [18:0] Wgt_8_101, // sfix19_En18 
  input [18:0] Wgt_8_102, // sfix19_En18 
  input [18:0] Wgt_8_103, // sfix19_En18 
  input [18:0] Wgt_8_104, // sfix19_En18 
  input [18:0] Wgt_8_105, // sfix19_En18 
  input [18:0] Wgt_8_106, // sfix19_En18 
  input [18:0] Wgt_8_107, // sfix19_En18 
  input [18:0] Wgt_8_108, // sfix19_En18 
  input [18:0] Wgt_8_109, // sfix19_En18 
  input [18:0] Wgt_8_110, // sfix19_En18 
  input [18:0] Wgt_8_111, // sfix19_En18 
  input [18:0] Wgt_8_112, // sfix19_En18 
  input [18:0] Wgt_8_113, // sfix19_En18 
  input [18:0] Wgt_8_114, // sfix19_En18 
  input [18:0] Wgt_8_115, // sfix19_En18 
  input [18:0] Wgt_8_116, // sfix19_En18 
  input [18:0] Wgt_8_117, // sfix19_En18 
  input [18:0] Wgt_8_118, // sfix19_En18 
  input [18:0] Wgt_8_119, // sfix19_En18 
  input [18:0] Wgt_8_120, // sfix19_En18 
  input [18:0] Wgt_8_121, // sfix19_En18 
  input [18:0] Wgt_8_122, // sfix19_En18 
  input [18:0] Wgt_8_123, // sfix19_En18 
  input [18:0] Wgt_8_124, // sfix19_En18 
  input [18:0] Wgt_8_125, // sfix19_En18 
  input [18:0] Wgt_8_126, // sfix19_En18 
  input [18:0] Wgt_8_127, // sfix19_En18 
  input [18:0] Wgt_8_128, // sfix19_En18 
  input [18:0] Wgt_8_129, // sfix19_En18 
  input [18:0] Wgt_8_130, // sfix19_En18 
  input [18:0] Wgt_8_131, // sfix19_En18 
  input [18:0] Wgt_8_132, // sfix19_En18 
  input [18:0] Wgt_8_133, // sfix19_En18 
  input [18:0] Wgt_8_134, // sfix19_En18 
  input [18:0] Wgt_8_135, // sfix19_En18 
  input [18:0] Wgt_8_136, // sfix19_En18 
  input [18:0] Wgt_8_137, // sfix19_En18 
  input [18:0] Wgt_8_138, // sfix19_En18 
  input [18:0] Wgt_8_139, // sfix19_En18 
  input [18:0] Wgt_8_140, // sfix19_En18 
  input [18:0] Wgt_8_141, // sfix19_En18 
  input [18:0] Wgt_8_142, // sfix19_En18 
  input [18:0] Wgt_8_143, // sfix19_En18 
  input [18:0] Wgt_8_144, // sfix19_En18 
  input [18:0] Wgt_8_145, // sfix19_En18 
  input [18:0] Wgt_8_146, // sfix19_En18 
  input [18:0] Wgt_8_147, // sfix19_En18 
  input [18:0] Wgt_8_148, // sfix19_En18 
  input [18:0] Wgt_8_149, // sfix19_En18 
  input [18:0] Wgt_8_150, // sfix19_En18 
  input [18:0] Wgt_8_151, // sfix19_En18 
  input [18:0] Wgt_8_152, // sfix19_En18 
  input [18:0] Wgt_8_153, // sfix19_En18 
  input [18:0] Wgt_8_154, // sfix19_En18 
  input [18:0] Wgt_8_155, // sfix19_En18 
  input [18:0] Wgt_8_156, // sfix19_En18 
  input [18:0] Wgt_8_157, // sfix19_En18 
  input [18:0] Wgt_8_158, // sfix19_En18 
  input [18:0] Wgt_8_159, // sfix19_En18 
  input [18:0] Wgt_8_160, // sfix19_En18 
  input [18:0] Wgt_8_161, // sfix19_En18 
  input [18:0] Wgt_8_162, // sfix19_En18 
  input [18:0] Wgt_8_163, // sfix19_En18 
  input [18:0] Wgt_8_164, // sfix19_En18 
  input [18:0] Wgt_8_165, // sfix19_En18 
  input [18:0] Wgt_8_166, // sfix19_En18 
  input [18:0] Wgt_8_167, // sfix19_En18 
  input [18:0] Wgt_8_168, // sfix19_En18 
  input [18:0] Wgt_8_169, // sfix19_En18 
  input [18:0] Wgt_8_170, // sfix19_En18 
  input [18:0] Wgt_8_171, // sfix19_En18 
  input [18:0] Wgt_8_172, // sfix19_En18 
  input [18:0] Wgt_8_173, // sfix19_En18 
  input [18:0] Wgt_8_174, // sfix19_En18 
  input [18:0] Wgt_8_175, // sfix19_En18 
  input [18:0] Wgt_8_176, // sfix19_En18 
  input [18:0] Wgt_8_177, // sfix19_En18 
  input [18:0] Wgt_8_178, // sfix19_En18 
  input [18:0] Wgt_8_179, // sfix19_En18 
  input [18:0] Wgt_8_180, // sfix19_En18 
  input [18:0] Wgt_8_181, // sfix19_En18 
  input [18:0] Wgt_8_182, // sfix19_En18 
  input [18:0] Wgt_8_183, // sfix19_En18 
  input [18:0] Wgt_8_184, // sfix19_En18 
  input [18:0] Wgt_8_185, // sfix19_En18 
  input [18:0] Wgt_8_186, // sfix19_En18 
  input [18:0] Wgt_8_187, // sfix19_En18 
  input [18:0] Wgt_8_188, // sfix19_En18 
  input [18:0] Wgt_8_189, // sfix19_En18 
  input [18:0] Wgt_8_190, // sfix19_En18 
  input [18:0] Wgt_8_191, // sfix19_En18 
  input [18:0] Wgt_8_192, // sfix19_En18 
  input [18:0] Wgt_8_193, // sfix19_En18 
  input [18:0] Wgt_8_194, // sfix19_En18 
  input [18:0] Wgt_8_195, // sfix19_En18 
  input [18:0] Wgt_8_196, // sfix19_En18 
  input [18:0] Wgt_8_197, // sfix19_En18 
  input [18:0] Wgt_8_198, // sfix19_En18 
  input [18:0] Wgt_8_199, // sfix19_En18 
  input [18:0] Wgt_8_200, // sfix19_En18 
  input [18:0] Wgt_8_201, // sfix19_En18 
  input [18:0] Wgt_8_202, // sfix19_En18 
  input [18:0] Wgt_8_203, // sfix19_En18 
  input [18:0] Wgt_8_204, // sfix19_En18 
  input [18:0] Wgt_8_205, // sfix19_En18 
  input [18:0] Wgt_8_206, // sfix19_En18 
  input [18:0] Wgt_8_207, // sfix19_En18 
  input [18:0] Wgt_8_208, // sfix19_En18 
  input [18:0] Wgt_8_209, // sfix19_En18 
  input [18:0] Wgt_8_210, // sfix19_En18 
  input [18:0] Wgt_8_211, // sfix19_En18 
  input [18:0] Wgt_8_212, // sfix19_En18 
  input [18:0] Wgt_8_213, // sfix19_En18 
  input [18:0] Wgt_8_214, // sfix19_En18 
  input [18:0] Wgt_8_215, // sfix19_En18 
  input [18:0] Wgt_8_216, // sfix19_En18 
  input [18:0] Wgt_8_217, // sfix19_En18 
  input [18:0] Wgt_8_218, // sfix19_En18 
  input [18:0] Wgt_8_219, // sfix19_En18 
  input [18:0] Wgt_8_220, // sfix19_En18 
  input [18:0] Wgt_8_221, // sfix19_En18 
  input [18:0] Wgt_8_222, // sfix19_En18 
  input [18:0] Wgt_8_223, // sfix19_En18 
  input [18:0] Wgt_8_224, // sfix19_En18 
  input [18:0] Wgt_8_225, // sfix19_En18 
  input [18:0] Wgt_8_226, // sfix19_En18 
  input [18:0] Wgt_8_227, // sfix19_En18 
  input [18:0] Wgt_8_228, // sfix19_En18 
  input [18:0] Wgt_8_229, // sfix19_En18 
  input [18:0] Wgt_8_230, // sfix19_En18 
  input [18:0] Wgt_8_231, // sfix19_En18 
  input [18:0] Wgt_8_232, // sfix19_En18 
  input [18:0] Wgt_8_233, // sfix19_En18 
  input [18:0] Wgt_8_234, // sfix19_En18 
  input [18:0] Wgt_8_235, // sfix19_En18 
  input [18:0] Wgt_8_236, // sfix19_En18 
  input [18:0] Wgt_8_237, // sfix19_En18 
  input [18:0] Wgt_8_238, // sfix19_En18 
  input [18:0] Wgt_8_239, // sfix19_En18 
  input [18:0] Wgt_8_240, // sfix19_En18 
  input [18:0] Wgt_8_241, // sfix19_En18 
  input [18:0] Wgt_8_242, // sfix19_En18 
  input [18:0] Wgt_8_243, // sfix19_En18 
  input [18:0] Wgt_8_244, // sfix19_En18 
  input [18:0] Wgt_8_245, // sfix19_En18 
  input [18:0] Wgt_8_246, // sfix19_En18 
  input [18:0] Wgt_8_247, // sfix19_En18 
  input [18:0] Wgt_8_248, // sfix19_En18 
  input [18:0] Wgt_8_249, // sfix19_En18 
  input [18:0] Wgt_8_250, // sfix19_En18 
  input [18:0] Wgt_8_251, // sfix19_En18 
  input [18:0] Wgt_8_252, // sfix19_En18 
  input [18:0] Wgt_8_253, // sfix19_En18 
  input [18:0] Wgt_8_254, // sfix19_En18 
  input [18:0] Wgt_8_255, // sfix19_En18 
  input [18:0] Wgt_8_256, // sfix19_En18 
  input [18:0] Wgt_8_257, // sfix19_En18 
  input [18:0] Wgt_8_258, // sfix19_En18 
  input [18:0] Wgt_8_259, // sfix19_En18 
  input [18:0] Wgt_8_260, // sfix19_En18 
  input [18:0] Wgt_8_261, // sfix19_En18 
  input [18:0] Wgt_8_262, // sfix19_En18 
  input [18:0] Wgt_8_263, // sfix19_En18 
  input [18:0] Wgt_8_264, // sfix19_En18 
  input [18:0] Wgt_8_265, // sfix19_En18 
  input [18:0] Wgt_8_266, // sfix19_En18 
  input [18:0] Wgt_8_267, // sfix19_En18 
  input [18:0] Wgt_8_268, // sfix19_En18 
  input [18:0] Wgt_8_269, // sfix19_En18 
  input [18:0] Wgt_8_270, // sfix19_En18 
  input [18:0] Wgt_8_271, // sfix19_En18 
  input [18:0] Wgt_8_272, // sfix19_En18 
  input [18:0] Wgt_8_273, // sfix19_En18 
  input [18:0] Wgt_8_274, // sfix19_En18 
  input [18:0] Wgt_8_275, // sfix19_En18 
  input [18:0] Wgt_8_276, // sfix19_En18 
  input [18:0] Wgt_8_277, // sfix19_En18 
  input [18:0] Wgt_8_278, // sfix19_En18 
  input [18:0] Wgt_8_279, // sfix19_En18 
  input [18:0] Wgt_8_280, // sfix19_En18 
  input [18:0] Wgt_8_281, // sfix19_En18 
  input [18:0] Wgt_8_282, // sfix19_En18 
  input [18:0] Wgt_8_283, // sfix19_En18 
  input [18:0] Wgt_8_284, // sfix19_En18 
  input [18:0] Wgt_8_285, // sfix19_En18 
  input [18:0] Wgt_8_286, // sfix19_En18 
  input [18:0] Wgt_8_287, // sfix19_En18 
  input [18:0] Wgt_8_288, // sfix19_En18 
  input [18:0] Wgt_8_289, // sfix19_En18 
  input [18:0] Wgt_8_290, // sfix19_En18 
  input [18:0] Wgt_8_291, // sfix19_En18 
  input [18:0] Wgt_8_292, // sfix19_En18 
  input [18:0] Wgt_8_293, // sfix19_En18 
  input [18:0] Wgt_8_294, // sfix19_En18 
  input [18:0] Wgt_8_295, // sfix19_En18 
  input [18:0] Wgt_8_296, // sfix19_En18 
  input [18:0] Wgt_8_297, // sfix19_En18 
  input [18:0] Wgt_8_298, // sfix19_En18 
  input [18:0] Wgt_8_299, // sfix19_En18 
  input [18:0] Wgt_8_300, // sfix19_En18 
  input [18:0] Wgt_8_301, // sfix19_En18 
  input [18:0] Wgt_8_302, // sfix19_En18 
  input [18:0] Wgt_8_303, // sfix19_En18 
  input [18:0] Wgt_8_304, // sfix19_En18 
  input [18:0] Wgt_8_305, // sfix19_En18 
  input [18:0] Wgt_8_306, // sfix19_En18 
  input [18:0] Wgt_8_307, // sfix19_En18 
  input [18:0] Wgt_8_308, // sfix19_En18 
  input [18:0] Wgt_8_309, // sfix19_En18 
  input [18:0] Wgt_8_310, // sfix19_En18 
  input [18:0] Wgt_8_311, // sfix19_En18 
  input [18:0] Wgt_8_312, // sfix19_En18 
  input [18:0] Wgt_8_313, // sfix19_En18 
  input [18:0] Wgt_8_314, // sfix19_En18 
  input [18:0] Wgt_8_315, // sfix19_En18 
  input [18:0] Wgt_8_316, // sfix19_En18 
  input [18:0] Wgt_8_317, // sfix19_En18 
  input [18:0] Wgt_8_318, // sfix19_En18 
  input [18:0] Wgt_8_319, // sfix19_En18 
  input [18:0] Wgt_8_320, // sfix19_En18 
  input [18:0] Wgt_8_321, // sfix19_En18 
  input [18:0] Wgt_8_322, // sfix19_En18 
  input [18:0] Wgt_8_323, // sfix19_En18 
  input [18:0] Wgt_8_324, // sfix19_En18 
  input [18:0] Wgt_8_325, // sfix19_En18 
  input [18:0] Wgt_8_326, // sfix19_En18 
  input [18:0] Wgt_8_327, // sfix19_En18 
  input [18:0] Wgt_8_328, // sfix19_En18 
  input [18:0] Wgt_8_329, // sfix19_En18 
  input [18:0] Wgt_8_330, // sfix19_En18 
  input [18:0] Wgt_8_331, // sfix19_En18 
  input [18:0] Wgt_8_332, // sfix19_En18 
  input [18:0] Wgt_8_333, // sfix19_En18 
  input [18:0] Wgt_8_334, // sfix19_En18 
  input [18:0] Wgt_8_335, // sfix19_En18 
  input [18:0] Wgt_8_336, // sfix19_En18 
  input [18:0] Wgt_8_337, // sfix19_En18 
  input [18:0] Wgt_8_338, // sfix19_En18 
  input [18:0] Wgt_8_339, // sfix19_En18 
  input [18:0] Wgt_8_340, // sfix19_En18 
  input [18:0] Wgt_8_341, // sfix19_En18 
  input [18:0] Wgt_8_342, // sfix19_En18 
  input [18:0] Wgt_8_343, // sfix19_En18 
  input [18:0] Wgt_8_344, // sfix19_En18 
  input [18:0] Wgt_8_345, // sfix19_En18 
  input [18:0] Wgt_8_346, // sfix19_En18 
  input [18:0] Wgt_8_347, // sfix19_En18 
  input [18:0] Wgt_8_348, // sfix19_En18 
  input [18:0] Wgt_8_349, // sfix19_En18 
  input [18:0] Wgt_8_350, // sfix19_En18 
  input [18:0] Wgt_8_351, // sfix19_En18 
  input [18:0] Wgt_8_352, // sfix19_En18 
  input [18:0] Wgt_8_353, // sfix19_En18 
  input [18:0] Wgt_8_354, // sfix19_En18 
  input [18:0] Wgt_8_355, // sfix19_En18 
  input [18:0] Wgt_8_356, // sfix19_En18 
  input [18:0] Wgt_8_357, // sfix19_En18 
  input [18:0] Wgt_8_358, // sfix19_En18 
  input [18:0] Wgt_8_359, // sfix19_En18 
  input [18:0] Wgt_8_360, // sfix19_En18 
  input [18:0] Wgt_8_361, // sfix19_En18 
  input [18:0] Wgt_8_362, // sfix19_En18 
  input [18:0] Wgt_8_363, // sfix19_En18 
  input [18:0] Wgt_8_364, // sfix19_En18 
  input [18:0] Wgt_8_365, // sfix19_En18 
  input [18:0] Wgt_8_366, // sfix19_En18 
  input [18:0] Wgt_8_367, // sfix19_En18 
  input [18:0] Wgt_8_368, // sfix19_En18 
  input [18:0] Wgt_8_369, // sfix19_En18 
  input [18:0] Wgt_8_370, // sfix19_En18 
  input [18:0] Wgt_8_371, // sfix19_En18 
  input [18:0] Wgt_8_372, // sfix19_En18 
  input [18:0] Wgt_8_373, // sfix19_En18 
  input [18:0] Wgt_8_374, // sfix19_En18 
  input [18:0] Wgt_8_375, // sfix19_En18 
  input [18:0] Wgt_8_376, // sfix19_En18 
  input [18:0] Wgt_8_377, // sfix19_En18 
  input [18:0] Wgt_8_378, // sfix19_En18 
  input [18:0] Wgt_8_379, // sfix19_En18 
  input [18:0] Wgt_8_380, // sfix19_En18 
  input [18:0] Wgt_8_381, // sfix19_En18 
  input [18:0] Wgt_8_382, // sfix19_En18 
  input [18:0] Wgt_8_383, // sfix19_En18 
  input [18:0] Wgt_8_384, // sfix19_En18 
  input [18:0] Wgt_8_385, // sfix19_En18 
  input [18:0] Wgt_8_386, // sfix19_En18 
  input [18:0] Wgt_8_387, // sfix19_En18 
  input [18:0] Wgt_8_388, // sfix19_En18 
  input [18:0] Wgt_8_389, // sfix19_En18 
  input [18:0] Wgt_8_390, // sfix19_En18 
  input [18:0] Wgt_8_391, // sfix19_En18 
  input [18:0] Wgt_8_392, // sfix19_En18 
  input [18:0] Wgt_8_393, // sfix19_En18 
  input [18:0] Wgt_8_394, // sfix19_En18 
  input [18:0] Wgt_8_395, // sfix19_En18 
  input [18:0] Wgt_8_396, // sfix19_En18 
  input [18:0] Wgt_8_397, // sfix19_En18 
  input [18:0] Wgt_8_398, // sfix19_En18 
  input [18:0] Wgt_8_399, // sfix19_En18 
  input [18:0] Wgt_8_400, // sfix19_En18 
  input [18:0] Wgt_8_401, // sfix19_En18 
  input [18:0] Wgt_8_402, // sfix19_En18 
  input [18:0] Wgt_8_403, // sfix19_En18 
  input [18:0] Wgt_8_404, // sfix19_En18 
  input [18:0] Wgt_8_405, // sfix19_En18 
  input [18:0] Wgt_8_406, // sfix19_En18 
  input [18:0] Wgt_8_407, // sfix19_En18 
  input [18:0] Wgt_8_408, // sfix19_En18 
  input [18:0] Wgt_8_409, // sfix19_En18 
  input [18:0] Wgt_8_410, // sfix19_En18 
  input [18:0] Wgt_8_411, // sfix19_En18 
  input [18:0] Wgt_8_412, // sfix19_En18 
  input [18:0] Wgt_8_413, // sfix19_En18 
  input [18:0] Wgt_8_414, // sfix19_En18 
  input [18:0] Wgt_8_415, // sfix19_En18 
  input [18:0] Wgt_8_416, // sfix19_En18 
  input [18:0] Wgt_8_417, // sfix19_En18 
  input [18:0] Wgt_8_418, // sfix19_En18 
  input [18:0] Wgt_8_419, // sfix19_En18 
  input [18:0] Wgt_8_420, // sfix19_En18 
  input [18:0] Wgt_8_421, // sfix19_En18 
  input [18:0] Wgt_8_422, // sfix19_En18 
  input [18:0] Wgt_8_423, // sfix19_En18 
  input [18:0] Wgt_8_424, // sfix19_En18 
  input [18:0] Wgt_8_425, // sfix19_En18 
  input [18:0] Wgt_8_426, // sfix19_En18 
  input [18:0] Wgt_8_427, // sfix19_En18 
  input [18:0] Wgt_8_428, // sfix19_En18 
  input [18:0] Wgt_8_429, // sfix19_En18 
  input [18:0] Wgt_8_430, // sfix19_En18 
  input [18:0] Wgt_8_431, // sfix19_En18 
  input [18:0] Wgt_8_432, // sfix19_En18 
  input [18:0] Wgt_8_433, // sfix19_En18 
  input [18:0] Wgt_8_434, // sfix19_En18 
  input [18:0] Wgt_8_435, // sfix19_En18 
  input [18:0] Wgt_8_436, // sfix19_En18 
  input [18:0] Wgt_8_437, // sfix19_En18 
  input [18:0] Wgt_8_438, // sfix19_En18 
  input [18:0] Wgt_8_439, // sfix19_En18 
  input [18:0] Wgt_8_440, // sfix19_En18 
  input [18:0] Wgt_8_441, // sfix19_En18 
  input [18:0] Wgt_8_442, // sfix19_En18 
  input [18:0] Wgt_8_443, // sfix19_En18 
  input [18:0] Wgt_8_444, // sfix19_En18 
  input [18:0] Wgt_8_445, // sfix19_En18 
  input [18:0] Wgt_8_446, // sfix19_En18 
  input [18:0] Wgt_8_447, // sfix19_En18 
  input [18:0] Wgt_8_448, // sfix19_En18 
  input [18:0] Wgt_8_449, // sfix19_En18 
  input [18:0] Wgt_8_450, // sfix19_En18 
  input [18:0] Wgt_8_451, // sfix19_En18 
  input [18:0] Wgt_8_452, // sfix19_En18 
  input [18:0] Wgt_8_453, // sfix19_En18 
  input [18:0] Wgt_8_454, // sfix19_En18 
  input [18:0] Wgt_8_455, // sfix19_En18 
  input [18:0] Wgt_8_456, // sfix19_En18 
  input [18:0] Wgt_8_457, // sfix19_En18 
  input [18:0] Wgt_8_458, // sfix19_En18 
  input [18:0] Wgt_8_459, // sfix19_En18 
  input [18:0] Wgt_8_460, // sfix19_En18 
  input [18:0] Wgt_8_461, // sfix19_En18 
  input [18:0] Wgt_8_462, // sfix19_En18 
  input [18:0] Wgt_8_463, // sfix19_En18 
  input [18:0] Wgt_8_464, // sfix19_En18 
  input [18:0] Wgt_8_465, // sfix19_En18 
  input [18:0] Wgt_8_466, // sfix19_En18 
  input [18:0] Wgt_8_467, // sfix19_En18 
  input [18:0] Wgt_8_468, // sfix19_En18 
  input [18:0] Wgt_8_469, // sfix19_En18 
  input [18:0] Wgt_8_470, // sfix19_En18 
  input [18:0] Wgt_8_471, // sfix19_En18 
  input [18:0] Wgt_8_472, // sfix19_En18 
  input [18:0] Wgt_8_473, // sfix19_En18 
  input [18:0] Wgt_8_474, // sfix19_En18 
  input [18:0] Wgt_8_475, // sfix19_En18 
  input [18:0] Wgt_8_476, // sfix19_En18 
  input [18:0] Wgt_8_477, // sfix19_En18 
  input [18:0] Wgt_8_478, // sfix19_En18 
  input [18:0] Wgt_8_479, // sfix19_En18 
  input [18:0] Wgt_8_480, // sfix19_En18 
  input [18:0] Wgt_8_481, // sfix19_En18 
  input [18:0] Wgt_8_482, // sfix19_En18 
  input [18:0] Wgt_8_483, // sfix19_En18 
  input [18:0] Wgt_8_484, // sfix19_En18 
  input [18:0] Wgt_8_485, // sfix19_En18 
  input [18:0] Wgt_8_486, // sfix19_En18 
  input [18:0] Wgt_8_487, // sfix19_En18 
  input [18:0] Wgt_8_488, // sfix19_En18 
  input [18:0] Wgt_8_489, // sfix19_En18 
  input [18:0] Wgt_8_490, // sfix19_En18 
  input [18:0] Wgt_8_491, // sfix19_En18 
  input [18:0] Wgt_8_492, // sfix19_En18 
  input [18:0] Wgt_8_493, // sfix19_En18 
  input [18:0] Wgt_8_494, // sfix19_En18 
  input [18:0] Wgt_8_495, // sfix19_En18 
  input [18:0] Wgt_8_496, // sfix19_En18 
  input [18:0] Wgt_8_497, // sfix19_En18 
  input [18:0] Wgt_8_498, // sfix19_En18 
  input [18:0] Wgt_8_499, // sfix19_En18 
  input [18:0] Wgt_8_500, // sfix19_En18 
  input [18:0] Wgt_8_501, // sfix19_En18 
  input [18:0] Wgt_8_502, // sfix19_En18 
  input [18:0] Wgt_8_503, // sfix19_En18 
  input [18:0] Wgt_8_504, // sfix19_En18 
  input [18:0] Wgt_8_505, // sfix19_En18 
  input [18:0] Wgt_8_506, // sfix19_En18 
  input [18:0] Wgt_8_507, // sfix19_En18 
  input [18:0] Wgt_8_508, // sfix19_En18 
  input [18:0] Wgt_8_509, // sfix19_En18 
  input [18:0] Wgt_8_510, // sfix19_En18 
  input [18:0] Wgt_8_511, // sfix19_En18 
  input [18:0] Wgt_8_512, // sfix19_En18 
  input [18:0] Wgt_8_513, // sfix19_En18 
  input [18:0] Wgt_8_514, // sfix19_En18 
  input [18:0] Wgt_8_515, // sfix19_En18 
  input [18:0] Wgt_8_516, // sfix19_En18 
  input [18:0] Wgt_8_517, // sfix19_En18 
  input [18:0] Wgt_8_518, // sfix19_En18 
  input [18:0] Wgt_8_519, // sfix19_En18 
  input [18:0] Wgt_8_520, // sfix19_En18 
  input [18:0] Wgt_8_521, // sfix19_En18 
  input [18:0] Wgt_8_522, // sfix19_En18 
  input [18:0] Wgt_8_523, // sfix19_En18 
  input [18:0] Wgt_8_524, // sfix19_En18 
  input [18:0] Wgt_8_525, // sfix19_En18 
  input [18:0] Wgt_8_526, // sfix19_En18 
  input [18:0] Wgt_8_527, // sfix19_En18 
  input [18:0] Wgt_8_528, // sfix19_En18 
  input [18:0] Wgt_8_529, // sfix19_En18 
  input [18:0] Wgt_8_530, // sfix19_En18 
  input [18:0] Wgt_8_531, // sfix19_En18 
  input [18:0] Wgt_8_532, // sfix19_En18 
  input [18:0] Wgt_8_533, // sfix19_En18 
  input [18:0] Wgt_8_534, // sfix19_En18 
  input [18:0] Wgt_8_535, // sfix19_En18 
  input [18:0] Wgt_8_536, // sfix19_En18 
  input [18:0] Wgt_8_537, // sfix19_En18 
  input [18:0] Wgt_8_538, // sfix19_En18 
  input [18:0] Wgt_8_539, // sfix19_En18 
  input [18:0] Wgt_8_540, // sfix19_En18 
  input [18:0] Wgt_8_541, // sfix19_En18 
  input [18:0] Wgt_8_542, // sfix19_En18 
  input [18:0] Wgt_8_543, // sfix19_En18 
  input [18:0] Wgt_8_544, // sfix19_En18 
  input [18:0] Wgt_8_545, // sfix19_En18 
  input [18:0] Wgt_8_546, // sfix19_En18 
  input [18:0] Wgt_8_547, // sfix19_En18 
  input [18:0] Wgt_8_548, // sfix19_En18 
  input [18:0] Wgt_8_549, // sfix19_En18 
  input [18:0] Wgt_8_550, // sfix19_En18 
  input [18:0] Wgt_8_551, // sfix19_En18 
  input [18:0] Wgt_8_552, // sfix19_En18 
  input [18:0] Wgt_8_553, // sfix19_En18 
  input [18:0] Wgt_8_554, // sfix19_En18 
  input [18:0] Wgt_8_555, // sfix19_En18 
  input [18:0] Wgt_8_556, // sfix19_En18 
  input [18:0] Wgt_8_557, // sfix19_En18 
  input [18:0] Wgt_8_558, // sfix19_En18 
  input [18:0] Wgt_8_559, // sfix19_En18 
  input [18:0] Wgt_8_560, // sfix19_En18 
  input [18:0] Wgt_8_561, // sfix19_En18 
  input [18:0] Wgt_8_562, // sfix19_En18 
  input [18:0] Wgt_8_563, // sfix19_En18 
  input [18:0] Wgt_8_564, // sfix19_En18 
  input [18:0] Wgt_8_565, // sfix19_En18 
  input [18:0] Wgt_8_566, // sfix19_En18 
  input [18:0] Wgt_8_567, // sfix19_En18 
  input [18:0] Wgt_8_568, // sfix19_En18 
  input [18:0] Wgt_8_569, // sfix19_En18 
  input [18:0] Wgt_8_570, // sfix19_En18 
  input [18:0] Wgt_8_571, // sfix19_En18 
  input [18:0] Wgt_8_572, // sfix19_En18 
  input [18:0] Wgt_8_573, // sfix19_En18 
  input [18:0] Wgt_8_574, // sfix19_En18 
  input [18:0] Wgt_8_575, // sfix19_En18 
  input [18:0] Wgt_8_576, // sfix19_En18 
  input [18:0] Wgt_8_577, // sfix19_En18 
  input [18:0] Wgt_8_578, // sfix19_En18 
  input [18:0] Wgt_8_579, // sfix19_En18 
  input [18:0] Wgt_8_580, // sfix19_En18 
  input [18:0] Wgt_8_581, // sfix19_En18 
  input [18:0] Wgt_8_582, // sfix19_En18 
  input [18:0] Wgt_8_583, // sfix19_En18 
  input [18:0] Wgt_8_584, // sfix19_En18 
  input [18:0] Wgt_8_585, // sfix19_En18 
  input [18:0] Wgt_8_586, // sfix19_En18 
  input [18:0] Wgt_8_587, // sfix19_En18 
  input [18:0] Wgt_8_588, // sfix19_En18 
  input [18:0] Wgt_8_589, // sfix19_En18 
  input [18:0] Wgt_8_590, // sfix19_En18 
  input [18:0] Wgt_8_591, // sfix19_En18 
  input [18:0] Wgt_8_592, // sfix19_En18 
  input [18:0] Wgt_8_593, // sfix19_En18 
  input [18:0] Wgt_8_594, // sfix19_En18 
  input [18:0] Wgt_8_595, // sfix19_En18 
  input [18:0] Wgt_8_596, // sfix19_En18 
  input [18:0] Wgt_8_597, // sfix19_En18 
  input [18:0] Wgt_8_598, // sfix19_En18 
  input [18:0] Wgt_8_599, // sfix19_En18 
  input [18:0] Wgt_8_600, // sfix19_En18 
  input [18:0] Wgt_8_601, // sfix19_En18 
  input [18:0] Wgt_8_602, // sfix19_En18 
  input [18:0] Wgt_8_603, // sfix19_En18 
  input [18:0] Wgt_8_604, // sfix19_En18 
  input [18:0] Wgt_8_605, // sfix19_En18 
  input [18:0] Wgt_8_606, // sfix19_En18 
  input [18:0] Wgt_8_607, // sfix19_En18 
  input [18:0] Wgt_8_608, // sfix19_En18 
  input [18:0] Wgt_8_609, // sfix19_En18 
  input [18:0] Wgt_8_610, // sfix19_En18 
  input [18:0] Wgt_8_611, // sfix19_En18 
  input [18:0] Wgt_8_612, // sfix19_En18 
  input [18:0] Wgt_8_613, // sfix19_En18 
  input [18:0] Wgt_8_614, // sfix19_En18 
  input [18:0] Wgt_8_615, // sfix19_En18 
  input [18:0] Wgt_8_616, // sfix19_En18 
  input [18:0] Wgt_8_617, // sfix19_En18 
  input [18:0] Wgt_8_618, // sfix19_En18 
  input [18:0] Wgt_8_619, // sfix19_En18 
  input [18:0] Wgt_8_620, // sfix19_En18 
  input [18:0] Wgt_8_621, // sfix19_En18 
  input [18:0] Wgt_8_622, // sfix19_En18 
  input [18:0] Wgt_8_623, // sfix19_En18 
  input [18:0] Wgt_8_624, // sfix19_En18 
  input [18:0] Wgt_8_625, // sfix19_En18 
  input [18:0] Wgt_8_626, // sfix19_En18 
  input [18:0] Wgt_8_627, // sfix19_En18 
  input [18:0] Wgt_8_628, // sfix19_En18 
  input [18:0] Wgt_8_629, // sfix19_En18 
  input [18:0] Wgt_8_630, // sfix19_En18 
  input [18:0] Wgt_8_631, // sfix19_En18 
  input [18:0] Wgt_8_632, // sfix19_En18 
  input [18:0] Wgt_8_633, // sfix19_En18 
  input [18:0] Wgt_8_634, // sfix19_En18 
  input [18:0] Wgt_8_635, // sfix19_En18 
  input [18:0] Wgt_8_636, // sfix19_En18 
  input [18:0] Wgt_8_637, // sfix19_En18 
  input [18:0] Wgt_8_638, // sfix19_En18 
  input [18:0] Wgt_8_639, // sfix19_En18 
  input [18:0] Wgt_8_640, // sfix19_En18 
  input [18:0] Wgt_8_641, // sfix19_En18 
  input [18:0] Wgt_8_642, // sfix19_En18 
  input [18:0] Wgt_8_643, // sfix19_En18 
  input [18:0] Wgt_8_644, // sfix19_En18 
  input [18:0] Wgt_8_645, // sfix19_En18 
  input [18:0] Wgt_8_646, // sfix19_En18 
  input [18:0] Wgt_8_647, // sfix19_En18 
  input [18:0] Wgt_8_648, // sfix19_En18 
  input [18:0] Wgt_8_649, // sfix19_En18 
  input [18:0] Wgt_8_650, // sfix19_En18 
  input [18:0] Wgt_8_651, // sfix19_En18 
  input [18:0] Wgt_8_652, // sfix19_En18 
  input [18:0] Wgt_8_653, // sfix19_En18 
  input [18:0] Wgt_8_654, // sfix19_En18 
  input [18:0] Wgt_8_655, // sfix19_En18 
  input [18:0] Wgt_8_656, // sfix19_En18 
  input [18:0] Wgt_8_657, // sfix19_En18 
  input [18:0] Wgt_8_658, // sfix19_En18 
  input [18:0] Wgt_8_659, // sfix19_En18 
  input [18:0] Wgt_8_660, // sfix19_En18 
  input [18:0] Wgt_8_661, // sfix19_En18 
  input [18:0] Wgt_8_662, // sfix19_En18 
  input [18:0] Wgt_8_663, // sfix19_En18 
  input [18:0] Wgt_8_664, // sfix19_En18 
  input [18:0] Wgt_8_665, // sfix19_En18 
  input [18:0] Wgt_8_666, // sfix19_En18 
  input [18:0] Wgt_8_667, // sfix19_En18 
  input [18:0] Wgt_8_668, // sfix19_En18 
  input [18:0] Wgt_8_669, // sfix19_En18 
  input [18:0] Wgt_8_670, // sfix19_En18 
  input [18:0] Wgt_8_671, // sfix19_En18 
  input [18:0] Wgt_8_672, // sfix19_En18 
  input [18:0] Wgt_8_673, // sfix19_En18 
  input [18:0] Wgt_8_674, // sfix19_En18 
  input [18:0] Wgt_8_675, // sfix19_En18 
  input [18:0] Wgt_8_676, // sfix19_En18 
  input [18:0] Wgt_8_677, // sfix19_En18 
  input [18:0] Wgt_8_678, // sfix19_En18 
  input [18:0] Wgt_8_679, // sfix19_En18 
  input [18:0] Wgt_8_680, // sfix19_En18 
  input [18:0] Wgt_8_681, // sfix19_En18 
  input [18:0] Wgt_8_682, // sfix19_En18 
  input [18:0] Wgt_8_683, // sfix19_En18 
  input [18:0] Wgt_8_684, // sfix19_En18 
  input [18:0] Wgt_8_685, // sfix19_En18 
  input [18:0] Wgt_8_686, // sfix19_En18 
  input [18:0] Wgt_8_687, // sfix19_En18 
  input [18:0] Wgt_8_688, // sfix19_En18 
  input [18:0] Wgt_8_689, // sfix19_En18 
  input [18:0] Wgt_8_690, // sfix19_En18 
  input [18:0] Wgt_8_691, // sfix19_En18 
  input [18:0] Wgt_8_692, // sfix19_En18 
  input [18:0] Wgt_8_693, // sfix19_En18 
  input [18:0] Wgt_8_694, // sfix19_En18 
  input [18:0] Wgt_8_695, // sfix19_En18 
  input [18:0] Wgt_8_696, // sfix19_En18 
  input [18:0] Wgt_8_697, // sfix19_En18 
  input [18:0] Wgt_8_698, // sfix19_En18 
  input [18:0] Wgt_8_699, // sfix19_En18 
  input [18:0] Wgt_8_700, // sfix19_En18 
  input [18:0] Wgt_8_701, // sfix19_En18 
  input [18:0] Wgt_8_702, // sfix19_En18 
  input [18:0] Wgt_8_703, // sfix19_En18 
  input [18:0] Wgt_8_704, // sfix19_En18 
  input [18:0] Wgt_8_705, // sfix19_En18 
  input [18:0] Wgt_8_706, // sfix19_En18 
  input [18:0] Wgt_8_707, // sfix19_En18 
  input [18:0] Wgt_8_708, // sfix19_En18 
  input [18:0] Wgt_8_709, // sfix19_En18 
  input [18:0] Wgt_8_710, // sfix19_En18 
  input [18:0] Wgt_8_711, // sfix19_En18 
  input [18:0] Wgt_8_712, // sfix19_En18 
  input [18:0] Wgt_8_713, // sfix19_En18 
  input [18:0] Wgt_8_714, // sfix19_En18 
  input [18:0] Wgt_8_715, // sfix19_En18 
  input [18:0] Wgt_8_716, // sfix19_En18 
  input [18:0] Wgt_8_717, // sfix19_En18 
  input [18:0] Wgt_8_718, // sfix19_En18 
  input [18:0] Wgt_8_719, // sfix19_En18 
  input [18:0] Wgt_8_720, // sfix19_En18 
  input [18:0] Wgt_8_721, // sfix19_En18 
  input [18:0] Wgt_8_722, // sfix19_En18 
  input [18:0] Wgt_8_723, // sfix19_En18 
  input [18:0] Wgt_8_724, // sfix19_En18 
  input [18:0] Wgt_8_725, // sfix19_En18 
  input [18:0] Wgt_8_726, // sfix19_En18 
  input [18:0] Wgt_8_727, // sfix19_En18 
  input [18:0] Wgt_8_728, // sfix19_En18 
  input [18:0] Wgt_8_729, // sfix19_En18 
  input [18:0] Wgt_8_730, // sfix19_En18 
  input [18:0] Wgt_8_731, // sfix19_En18 
  input [18:0] Wgt_8_732, // sfix19_En18 
  input [18:0] Wgt_8_733, // sfix19_En18 
  input [18:0] Wgt_8_734, // sfix19_En18 
  input [18:0] Wgt_8_735, // sfix19_En18 
  input [18:0] Wgt_8_736, // sfix19_En18 
  input [18:0] Wgt_8_737, // sfix19_En18 
  input [18:0] Wgt_8_738, // sfix19_En18 
  input [18:0] Wgt_8_739, // sfix19_En18 
  input [18:0] Wgt_8_740, // sfix19_En18 
  input [18:0] Wgt_8_741, // sfix19_En18 
  input [18:0] Wgt_8_742, // sfix19_En18 
  input [18:0] Wgt_8_743, // sfix19_En18 
  input [18:0] Wgt_8_744, // sfix19_En18 
  input [18:0] Wgt_8_745, // sfix19_En18 
  input [18:0] Wgt_8_746, // sfix19_En18 
  input [18:0] Wgt_8_747, // sfix19_En18 
  input [18:0] Wgt_8_748, // sfix19_En18 
  input [18:0] Wgt_8_749, // sfix19_En18 
  input [18:0] Wgt_8_750, // sfix19_En18 
  input [18:0] Wgt_8_751, // sfix19_En18 
  input [18:0] Wgt_8_752, // sfix19_En18 
  input [18:0] Wgt_8_753, // sfix19_En18 
  input [18:0] Wgt_8_754, // sfix19_En18 
  input [18:0] Wgt_8_755, // sfix19_En18 
  input [18:0] Wgt_8_756, // sfix19_En18 
  input [18:0] Wgt_8_757, // sfix19_En18 
  input [18:0] Wgt_8_758, // sfix19_En18 
  input [18:0] Wgt_8_759, // sfix19_En18 
  input [18:0] Wgt_8_760, // sfix19_En18 
  input [18:0] Wgt_8_761, // sfix19_En18 
  input [18:0] Wgt_8_762, // sfix19_En18 
  input [18:0] Wgt_8_763, // sfix19_En18 
  input [18:0] Wgt_8_764, // sfix19_En18 
  input [18:0] Wgt_8_765, // sfix19_En18 
  input [18:0] Wgt_8_766, // sfix19_En18 
  input [18:0] Wgt_8_767, // sfix19_En18 
  input [18:0] Wgt_8_768, // sfix19_En18 
  input [18:0] Wgt_8_769, // sfix19_En18 
  input [18:0] Wgt_8_770, // sfix19_En18 
  input [18:0] Wgt_8_771, // sfix19_En18 
  input [18:0] Wgt_8_772, // sfix19_En18 
  input [18:0] Wgt_8_773, // sfix19_En18 
  input [18:0] Wgt_8_774, // sfix19_En18 
  input [18:0] Wgt_8_775, // sfix19_En18 
  input [18:0] Wgt_8_776, // sfix19_En18 
  input [18:0] Wgt_8_777, // sfix19_En18 
  input [18:0] Wgt_8_778, // sfix19_En18 
  input [18:0] Wgt_8_779, // sfix19_En18 
  input [18:0] Wgt_8_780, // sfix19_En18 
  input [18:0] Wgt_8_781, // sfix19_En18 
  input [18:0] Wgt_8_782, // sfix19_En18 
  input [18:0] Wgt_8_783, // sfix19_En18 
  input [18:0] Wgt_8_784, // sfix19_En18 
  input [18:0] Wgt_9_0, // sfix19_En18 
  input [18:0] Wgt_9_1, // sfix19_En18 
  input [18:0] Wgt_9_2, // sfix19_En18 
  input [18:0] Wgt_9_3, // sfix19_En18 
  input [18:0] Wgt_9_4, // sfix19_En18 
  input [18:0] Wgt_9_5, // sfix19_En18 
  input [18:0] Wgt_9_6, // sfix19_En18 
  input [18:0] Wgt_9_7, // sfix19_En18 
  input [18:0] Wgt_9_8, // sfix19_En18 
  input [18:0] Wgt_9_9, // sfix19_En18 
  input [18:0] Wgt_9_10, // sfix19_En18 
  input [18:0] Wgt_9_11, // sfix19_En18 
  input [18:0] Wgt_9_12, // sfix19_En18 
  input [18:0] Wgt_9_13, // sfix19_En18 
  input [18:0] Wgt_9_14, // sfix19_En18 
  input [18:0] Wgt_9_15, // sfix19_En18 
  input [18:0] Wgt_9_16, // sfix19_En18 
  input [18:0] Wgt_9_17, // sfix19_En18 
  input [18:0] Wgt_9_18, // sfix19_En18 
  input [18:0] Wgt_9_19, // sfix19_En18 
  input [18:0] Wgt_9_20, // sfix19_En18 
  input [18:0] Wgt_9_21, // sfix19_En18 
  input [18:0] Wgt_9_22, // sfix19_En18 
  input [18:0] Wgt_9_23, // sfix19_En18 
  input [18:0] Wgt_9_24, // sfix19_En18 
  input [18:0] Wgt_9_25, // sfix19_En18 
  input [18:0] Wgt_9_26, // sfix19_En18 
  input [18:0] Wgt_9_27, // sfix19_En18 
  input [18:0] Wgt_9_28, // sfix19_En18 
  input [18:0] Wgt_9_29, // sfix19_En18 
  input [18:0] Wgt_9_30, // sfix19_En18 
  input [18:0] Wgt_9_31, // sfix19_En18 
  input [18:0] Wgt_9_32, // sfix19_En18 
  input [18:0] Wgt_9_33, // sfix19_En18 
  input [18:0] Wgt_9_34, // sfix19_En18 
  input [18:0] Wgt_9_35, // sfix19_En18 
  input [18:0] Wgt_9_36, // sfix19_En18 
  input [18:0] Wgt_9_37, // sfix19_En18 
  input [18:0] Wgt_9_38, // sfix19_En18 
  input [18:0] Wgt_9_39, // sfix19_En18 
  input [18:0] Wgt_9_40, // sfix19_En18 
  input [18:0] Wgt_9_41, // sfix19_En18 
  input [18:0] Wgt_9_42, // sfix19_En18 
  input [18:0] Wgt_9_43, // sfix19_En18 
  input [18:0] Wgt_9_44, // sfix19_En18 
  input [18:0] Wgt_9_45, // sfix19_En18 
  input [18:0] Wgt_9_46, // sfix19_En18 
  input [18:0] Wgt_9_47, // sfix19_En18 
  input [18:0] Wgt_9_48, // sfix19_En18 
  input [18:0] Wgt_9_49, // sfix19_En18 
  input [18:0] Wgt_9_50, // sfix19_En18 
  input [18:0] Wgt_9_51, // sfix19_En18 
  input [18:0] Wgt_9_52, // sfix19_En18 
  input [18:0] Wgt_9_53, // sfix19_En18 
  input [18:0] Wgt_9_54, // sfix19_En18 
  input [18:0] Wgt_9_55, // sfix19_En18 
  input [18:0] Wgt_9_56, // sfix19_En18 
  input [18:0] Wgt_9_57, // sfix19_En18 
  input [18:0] Wgt_9_58, // sfix19_En18 
  input [18:0] Wgt_9_59, // sfix19_En18 
  input [18:0] Wgt_9_60, // sfix19_En18 
  input [18:0] Wgt_9_61, // sfix19_En18 
  input [18:0] Wgt_9_62, // sfix19_En18 
  input [18:0] Wgt_9_63, // sfix19_En18 
  input [18:0] Wgt_9_64, // sfix19_En18 
  input [18:0] Wgt_9_65, // sfix19_En18 
  input [18:0] Wgt_9_66, // sfix19_En18 
  input [18:0] Wgt_9_67, // sfix19_En18 
  input [18:0] Wgt_9_68, // sfix19_En18 
  input [18:0] Wgt_9_69, // sfix19_En18 
  input [18:0] Wgt_9_70, // sfix19_En18 
  input [18:0] Wgt_9_71, // sfix19_En18 
  input [18:0] Wgt_9_72, // sfix19_En18 
  input [18:0] Wgt_9_73, // sfix19_En18 
  input [18:0] Wgt_9_74, // sfix19_En18 
  input [18:0] Wgt_9_75, // sfix19_En18 
  input [18:0] Wgt_9_76, // sfix19_En18 
  input [18:0] Wgt_9_77, // sfix19_En18 
  input [18:0] Wgt_9_78, // sfix19_En18 
  input [18:0] Wgt_9_79, // sfix19_En18 
  input [18:0] Wgt_9_80, // sfix19_En18 
  input [18:0] Wgt_9_81, // sfix19_En18 
  input [18:0] Wgt_9_82, // sfix19_En18 
  input [18:0] Wgt_9_83, // sfix19_En18 
  input [18:0] Wgt_9_84, // sfix19_En18 
  input [18:0] Wgt_9_85, // sfix19_En18 
  input [18:0] Wgt_9_86, // sfix19_En18 
  input [18:0] Wgt_9_87, // sfix19_En18 
  input [18:0] Wgt_9_88, // sfix19_En18 
  input [18:0] Wgt_9_89, // sfix19_En18 
  input [18:0] Wgt_9_90, // sfix19_En18 
  input [18:0] Wgt_9_91, // sfix19_En18 
  input [18:0] Wgt_9_92, // sfix19_En18 
  input [18:0] Wgt_9_93, // sfix19_En18 
  input [18:0] Wgt_9_94, // sfix19_En18 
  input [18:0] Wgt_9_95, // sfix19_En18 
  input [18:0] Wgt_9_96, // sfix19_En18 
  input [18:0] Wgt_9_97, // sfix19_En18 
  input [18:0] Wgt_9_98, // sfix19_En18 
  input [18:0] Wgt_9_99, // sfix19_En18 
  input [18:0] Wgt_9_100, // sfix19_En18 
  input [18:0] Wgt_9_101, // sfix19_En18 
  input [18:0] Wgt_9_102, // sfix19_En18 
  input [18:0] Wgt_9_103, // sfix19_En18 
  input [18:0] Wgt_9_104, // sfix19_En18 
  input [18:0] Wgt_9_105, // sfix19_En18 
  input [18:0] Wgt_9_106, // sfix19_En18 
  input [18:0] Wgt_9_107, // sfix19_En18 
  input [18:0] Wgt_9_108, // sfix19_En18 
  input [18:0] Wgt_9_109, // sfix19_En18 
  input [18:0] Wgt_9_110, // sfix19_En18 
  input [18:0] Wgt_9_111, // sfix19_En18 
  input [18:0] Wgt_9_112, // sfix19_En18 
  input [18:0] Wgt_9_113, // sfix19_En18 
  input [18:0] Wgt_9_114, // sfix19_En18 
  input [18:0] Wgt_9_115, // sfix19_En18 
  input [18:0] Wgt_9_116, // sfix19_En18 
  input [18:0] Wgt_9_117, // sfix19_En18 
  input [18:0] Wgt_9_118, // sfix19_En18 
  input [18:0] Wgt_9_119, // sfix19_En18 
  input [18:0] Wgt_9_120, // sfix19_En18 
  input [18:0] Wgt_9_121, // sfix19_En18 
  input [18:0] Wgt_9_122, // sfix19_En18 
  input [18:0] Wgt_9_123, // sfix19_En18 
  input [18:0] Wgt_9_124, // sfix19_En18 
  input [18:0] Wgt_9_125, // sfix19_En18 
  input [18:0] Wgt_9_126, // sfix19_En18 
  input [18:0] Wgt_9_127, // sfix19_En18 
  input [18:0] Wgt_9_128, // sfix19_En18 
  input [18:0] Wgt_9_129, // sfix19_En18 
  input [18:0] Wgt_9_130, // sfix19_En18 
  input [18:0] Wgt_9_131, // sfix19_En18 
  input [18:0] Wgt_9_132, // sfix19_En18 
  input [18:0] Wgt_9_133, // sfix19_En18 
  input [18:0] Wgt_9_134, // sfix19_En18 
  input [18:0] Wgt_9_135, // sfix19_En18 
  input [18:0] Wgt_9_136, // sfix19_En18 
  input [18:0] Wgt_9_137, // sfix19_En18 
  input [18:0] Wgt_9_138, // sfix19_En18 
  input [18:0] Wgt_9_139, // sfix19_En18 
  input [18:0] Wgt_9_140, // sfix19_En18 
  input [18:0] Wgt_9_141, // sfix19_En18 
  input [18:0] Wgt_9_142, // sfix19_En18 
  input [18:0] Wgt_9_143, // sfix19_En18 
  input [18:0] Wgt_9_144, // sfix19_En18 
  input [18:0] Wgt_9_145, // sfix19_En18 
  input [18:0] Wgt_9_146, // sfix19_En18 
  input [18:0] Wgt_9_147, // sfix19_En18 
  input [18:0] Wgt_9_148, // sfix19_En18 
  input [18:0] Wgt_9_149, // sfix19_En18 
  input [18:0] Wgt_9_150, // sfix19_En18 
  input [18:0] Wgt_9_151, // sfix19_En18 
  input [18:0] Wgt_9_152, // sfix19_En18 
  input [18:0] Wgt_9_153, // sfix19_En18 
  input [18:0] Wgt_9_154, // sfix19_En18 
  input [18:0] Wgt_9_155, // sfix19_En18 
  input [18:0] Wgt_9_156, // sfix19_En18 
  input [18:0] Wgt_9_157, // sfix19_En18 
  input [18:0] Wgt_9_158, // sfix19_En18 
  input [18:0] Wgt_9_159, // sfix19_En18 
  input [18:0] Wgt_9_160, // sfix19_En18 
  input [18:0] Wgt_9_161, // sfix19_En18 
  input [18:0] Wgt_9_162, // sfix19_En18 
  input [18:0] Wgt_9_163, // sfix19_En18 
  input [18:0] Wgt_9_164, // sfix19_En18 
  input [18:0] Wgt_9_165, // sfix19_En18 
  input [18:0] Wgt_9_166, // sfix19_En18 
  input [18:0] Wgt_9_167, // sfix19_En18 
  input [18:0] Wgt_9_168, // sfix19_En18 
  input [18:0] Wgt_9_169, // sfix19_En18 
  input [18:0] Wgt_9_170, // sfix19_En18 
  input [18:0] Wgt_9_171, // sfix19_En18 
  input [18:0] Wgt_9_172, // sfix19_En18 
  input [18:0] Wgt_9_173, // sfix19_En18 
  input [18:0] Wgt_9_174, // sfix19_En18 
  input [18:0] Wgt_9_175, // sfix19_En18 
  input [18:0] Wgt_9_176, // sfix19_En18 
  input [18:0] Wgt_9_177, // sfix19_En18 
  input [18:0] Wgt_9_178, // sfix19_En18 
  input [18:0] Wgt_9_179, // sfix19_En18 
  input [18:0] Wgt_9_180, // sfix19_En18 
  input [18:0] Wgt_9_181, // sfix19_En18 
  input [18:0] Wgt_9_182, // sfix19_En18 
  input [18:0] Wgt_9_183, // sfix19_En18 
  input [18:0] Wgt_9_184, // sfix19_En18 
  input [18:0] Wgt_9_185, // sfix19_En18 
  input [18:0] Wgt_9_186, // sfix19_En18 
  input [18:0] Wgt_9_187, // sfix19_En18 
  input [18:0] Wgt_9_188, // sfix19_En18 
  input [18:0] Wgt_9_189, // sfix19_En18 
  input [18:0] Wgt_9_190, // sfix19_En18 
  input [18:0] Wgt_9_191, // sfix19_En18 
  input [18:0] Wgt_9_192, // sfix19_En18 
  input [18:0] Wgt_9_193, // sfix19_En18 
  input [18:0] Wgt_9_194, // sfix19_En18 
  input [18:0] Wgt_9_195, // sfix19_En18 
  input [18:0] Wgt_9_196, // sfix19_En18 
  input [18:0] Wgt_9_197, // sfix19_En18 
  input [18:0] Wgt_9_198, // sfix19_En18 
  input [18:0] Wgt_9_199, // sfix19_En18 
  input [18:0] Wgt_9_200, // sfix19_En18 
  input [18:0] Wgt_9_201, // sfix19_En18 
  input [18:0] Wgt_9_202, // sfix19_En18 
  input [18:0] Wgt_9_203, // sfix19_En18 
  input [18:0] Wgt_9_204, // sfix19_En18 
  input [18:0] Wgt_9_205, // sfix19_En18 
  input [18:0] Wgt_9_206, // sfix19_En18 
  input [18:0] Wgt_9_207, // sfix19_En18 
  input [18:0] Wgt_9_208, // sfix19_En18 
  input [18:0] Wgt_9_209, // sfix19_En18 
  input [18:0] Wgt_9_210, // sfix19_En18 
  input [18:0] Wgt_9_211, // sfix19_En18 
  input [18:0] Wgt_9_212, // sfix19_En18 
  input [18:0] Wgt_9_213, // sfix19_En18 
  input [18:0] Wgt_9_214, // sfix19_En18 
  input [18:0] Wgt_9_215, // sfix19_En18 
  input [18:0] Wgt_9_216, // sfix19_En18 
  input [18:0] Wgt_9_217, // sfix19_En18 
  input [18:0] Wgt_9_218, // sfix19_En18 
  input [18:0] Wgt_9_219, // sfix19_En18 
  input [18:0] Wgt_9_220, // sfix19_En18 
  input [18:0] Wgt_9_221, // sfix19_En18 
  input [18:0] Wgt_9_222, // sfix19_En18 
  input [18:0] Wgt_9_223, // sfix19_En18 
  input [18:0] Wgt_9_224, // sfix19_En18 
  input [18:0] Wgt_9_225, // sfix19_En18 
  input [18:0] Wgt_9_226, // sfix19_En18 
  input [18:0] Wgt_9_227, // sfix19_En18 
  input [18:0] Wgt_9_228, // sfix19_En18 
  input [18:0] Wgt_9_229, // sfix19_En18 
  input [18:0] Wgt_9_230, // sfix19_En18 
  input [18:0] Wgt_9_231, // sfix19_En18 
  input [18:0] Wgt_9_232, // sfix19_En18 
  input [18:0] Wgt_9_233, // sfix19_En18 
  input [18:0] Wgt_9_234, // sfix19_En18 
  input [18:0] Wgt_9_235, // sfix19_En18 
  input [18:0] Wgt_9_236, // sfix19_En18 
  input [18:0] Wgt_9_237, // sfix19_En18 
  input [18:0] Wgt_9_238, // sfix19_En18 
  input [18:0] Wgt_9_239, // sfix19_En18 
  input [18:0] Wgt_9_240, // sfix19_En18 
  input [18:0] Wgt_9_241, // sfix19_En18 
  input [18:0] Wgt_9_242, // sfix19_En18 
  input [18:0] Wgt_9_243, // sfix19_En18 
  input [18:0] Wgt_9_244, // sfix19_En18 
  input [18:0] Wgt_9_245, // sfix19_En18 
  input [18:0] Wgt_9_246, // sfix19_En18 
  input [18:0] Wgt_9_247, // sfix19_En18 
  input [18:0] Wgt_9_248, // sfix19_En18 
  input [18:0] Wgt_9_249, // sfix19_En18 
  input [18:0] Wgt_9_250, // sfix19_En18 
  input [18:0] Wgt_9_251, // sfix19_En18 
  input [18:0] Wgt_9_252, // sfix19_En18 
  input [18:0] Wgt_9_253, // sfix19_En18 
  input [18:0] Wgt_9_254, // sfix19_En18 
  input [18:0] Wgt_9_255, // sfix19_En18 
  input [18:0] Wgt_9_256, // sfix19_En18 
  input [18:0] Wgt_9_257, // sfix19_En18 
  input [18:0] Wgt_9_258, // sfix19_En18 
  input [18:0] Wgt_9_259, // sfix19_En18 
  input [18:0] Wgt_9_260, // sfix19_En18 
  input [18:0] Wgt_9_261, // sfix19_En18 
  input [18:0] Wgt_9_262, // sfix19_En18 
  input [18:0] Wgt_9_263, // sfix19_En18 
  input [18:0] Wgt_9_264, // sfix19_En18 
  input [18:0] Wgt_9_265, // sfix19_En18 
  input [18:0] Wgt_9_266, // sfix19_En18 
  input [18:0] Wgt_9_267, // sfix19_En18 
  input [18:0] Wgt_9_268, // sfix19_En18 
  input [18:0] Wgt_9_269, // sfix19_En18 
  input [18:0] Wgt_9_270, // sfix19_En18 
  input [18:0] Wgt_9_271, // sfix19_En18 
  input [18:0] Wgt_9_272, // sfix19_En18 
  input [18:0] Wgt_9_273, // sfix19_En18 
  input [18:0] Wgt_9_274, // sfix19_En18 
  input [18:0] Wgt_9_275, // sfix19_En18 
  input [18:0] Wgt_9_276, // sfix19_En18 
  input [18:0] Wgt_9_277, // sfix19_En18 
  input [18:0] Wgt_9_278, // sfix19_En18 
  input [18:0] Wgt_9_279, // sfix19_En18 
  input [18:0] Wgt_9_280, // sfix19_En18 
  input [18:0] Wgt_9_281, // sfix19_En18 
  input [18:0] Wgt_9_282, // sfix19_En18 
  input [18:0] Wgt_9_283, // sfix19_En18 
  input [18:0] Wgt_9_284, // sfix19_En18 
  input [18:0] Wgt_9_285, // sfix19_En18 
  input [18:0] Wgt_9_286, // sfix19_En18 
  input [18:0] Wgt_9_287, // sfix19_En18 
  input [18:0] Wgt_9_288, // sfix19_En18 
  input [18:0] Wgt_9_289, // sfix19_En18 
  input [18:0] Wgt_9_290, // sfix19_En18 
  input [18:0] Wgt_9_291, // sfix19_En18 
  input [18:0] Wgt_9_292, // sfix19_En18 
  input [18:0] Wgt_9_293, // sfix19_En18 
  input [18:0] Wgt_9_294, // sfix19_En18 
  input [18:0] Wgt_9_295, // sfix19_En18 
  input [18:0] Wgt_9_296, // sfix19_En18 
  input [18:0] Wgt_9_297, // sfix19_En18 
  input [18:0] Wgt_9_298, // sfix19_En18 
  input [18:0] Wgt_9_299, // sfix19_En18 
  input [18:0] Wgt_9_300, // sfix19_En18 
  input [18:0] Wgt_9_301, // sfix19_En18 
  input [18:0] Wgt_9_302, // sfix19_En18 
  input [18:0] Wgt_9_303, // sfix19_En18 
  input [18:0] Wgt_9_304, // sfix19_En18 
  input [18:0] Wgt_9_305, // sfix19_En18 
  input [18:0] Wgt_9_306, // sfix19_En18 
  input [18:0] Wgt_9_307, // sfix19_En18 
  input [18:0] Wgt_9_308, // sfix19_En18 
  input [18:0] Wgt_9_309, // sfix19_En18 
  input [18:0] Wgt_9_310, // sfix19_En18 
  input [18:0] Wgt_9_311, // sfix19_En18 
  input [18:0] Wgt_9_312, // sfix19_En18 
  input [18:0] Wgt_9_313, // sfix19_En18 
  input [18:0] Wgt_9_314, // sfix19_En18 
  input [18:0] Wgt_9_315, // sfix19_En18 
  input [18:0] Wgt_9_316, // sfix19_En18 
  input [18:0] Wgt_9_317, // sfix19_En18 
  input [18:0] Wgt_9_318, // sfix19_En18 
  input [18:0] Wgt_9_319, // sfix19_En18 
  input [18:0] Wgt_9_320, // sfix19_En18 
  input [18:0] Wgt_9_321, // sfix19_En18 
  input [18:0] Wgt_9_322, // sfix19_En18 
  input [18:0] Wgt_9_323, // sfix19_En18 
  input [18:0] Wgt_9_324, // sfix19_En18 
  input [18:0] Wgt_9_325, // sfix19_En18 
  input [18:0] Wgt_9_326, // sfix19_En18 
  input [18:0] Wgt_9_327, // sfix19_En18 
  input [18:0] Wgt_9_328, // sfix19_En18 
  input [18:0] Wgt_9_329, // sfix19_En18 
  input [18:0] Wgt_9_330, // sfix19_En18 
  input [18:0] Wgt_9_331, // sfix19_En18 
  input [18:0] Wgt_9_332, // sfix19_En18 
  input [18:0] Wgt_9_333, // sfix19_En18 
  input [18:0] Wgt_9_334, // sfix19_En18 
  input [18:0] Wgt_9_335, // sfix19_En18 
  input [18:0] Wgt_9_336, // sfix19_En18 
  input [18:0] Wgt_9_337, // sfix19_En18 
  input [18:0] Wgt_9_338, // sfix19_En18 
  input [18:0] Wgt_9_339, // sfix19_En18 
  input [18:0] Wgt_9_340, // sfix19_En18 
  input [18:0] Wgt_9_341, // sfix19_En18 
  input [18:0] Wgt_9_342, // sfix19_En18 
  input [18:0] Wgt_9_343, // sfix19_En18 
  input [18:0] Wgt_9_344, // sfix19_En18 
  input [18:0] Wgt_9_345, // sfix19_En18 
  input [18:0] Wgt_9_346, // sfix19_En18 
  input [18:0] Wgt_9_347, // sfix19_En18 
  input [18:0] Wgt_9_348, // sfix19_En18 
  input [18:0] Wgt_9_349, // sfix19_En18 
  input [18:0] Wgt_9_350, // sfix19_En18 
  input [18:0] Wgt_9_351, // sfix19_En18 
  input [18:0] Wgt_9_352, // sfix19_En18 
  input [18:0] Wgt_9_353, // sfix19_En18 
  input [18:0] Wgt_9_354, // sfix19_En18 
  input [18:0] Wgt_9_355, // sfix19_En18 
  input [18:0] Wgt_9_356, // sfix19_En18 
  input [18:0] Wgt_9_357, // sfix19_En18 
  input [18:0] Wgt_9_358, // sfix19_En18 
  input [18:0] Wgt_9_359, // sfix19_En18 
  input [18:0] Wgt_9_360, // sfix19_En18 
  input [18:0] Wgt_9_361, // sfix19_En18 
  input [18:0] Wgt_9_362, // sfix19_En18 
  input [18:0] Wgt_9_363, // sfix19_En18 
  input [18:0] Wgt_9_364, // sfix19_En18 
  input [18:0] Wgt_9_365, // sfix19_En18 
  input [18:0] Wgt_9_366, // sfix19_En18 
  input [18:0] Wgt_9_367, // sfix19_En18 
  input [18:0] Wgt_9_368, // sfix19_En18 
  input [18:0] Wgt_9_369, // sfix19_En18 
  input [18:0] Wgt_9_370, // sfix19_En18 
  input [18:0] Wgt_9_371, // sfix19_En18 
  input [18:0] Wgt_9_372, // sfix19_En18 
  input [18:0] Wgt_9_373, // sfix19_En18 
  input [18:0] Wgt_9_374, // sfix19_En18 
  input [18:0] Wgt_9_375, // sfix19_En18 
  input [18:0] Wgt_9_376, // sfix19_En18 
  input [18:0] Wgt_9_377, // sfix19_En18 
  input [18:0] Wgt_9_378, // sfix19_En18 
  input [18:0] Wgt_9_379, // sfix19_En18 
  input [18:0] Wgt_9_380, // sfix19_En18 
  input [18:0] Wgt_9_381, // sfix19_En18 
  input [18:0] Wgt_9_382, // sfix19_En18 
  input [18:0] Wgt_9_383, // sfix19_En18 
  input [18:0] Wgt_9_384, // sfix19_En18 
  input [18:0] Wgt_9_385, // sfix19_En18 
  input [18:0] Wgt_9_386, // sfix19_En18 
  input [18:0] Wgt_9_387, // sfix19_En18 
  input [18:0] Wgt_9_388, // sfix19_En18 
  input [18:0] Wgt_9_389, // sfix19_En18 
  input [18:0] Wgt_9_390, // sfix19_En18 
  input [18:0] Wgt_9_391, // sfix19_En18 
  input [18:0] Wgt_9_392, // sfix19_En18 
  input [18:0] Wgt_9_393, // sfix19_En18 
  input [18:0] Wgt_9_394, // sfix19_En18 
  input [18:0] Wgt_9_395, // sfix19_En18 
  input [18:0] Wgt_9_396, // sfix19_En18 
  input [18:0] Wgt_9_397, // sfix19_En18 
  input [18:0] Wgt_9_398, // sfix19_En18 
  input [18:0] Wgt_9_399, // sfix19_En18 
  input [18:0] Wgt_9_400, // sfix19_En18 
  input [18:0] Wgt_9_401, // sfix19_En18 
  input [18:0] Wgt_9_402, // sfix19_En18 
  input [18:0] Wgt_9_403, // sfix19_En18 
  input [18:0] Wgt_9_404, // sfix19_En18 
  input [18:0] Wgt_9_405, // sfix19_En18 
  input [18:0] Wgt_9_406, // sfix19_En18 
  input [18:0] Wgt_9_407, // sfix19_En18 
  input [18:0] Wgt_9_408, // sfix19_En18 
  input [18:0] Wgt_9_409, // sfix19_En18 
  input [18:0] Wgt_9_410, // sfix19_En18 
  input [18:0] Wgt_9_411, // sfix19_En18 
  input [18:0] Wgt_9_412, // sfix19_En18 
  input [18:0] Wgt_9_413, // sfix19_En18 
  input [18:0] Wgt_9_414, // sfix19_En18 
  input [18:0] Wgt_9_415, // sfix19_En18 
  input [18:0] Wgt_9_416, // sfix19_En18 
  input [18:0] Wgt_9_417, // sfix19_En18 
  input [18:0] Wgt_9_418, // sfix19_En18 
  input [18:0] Wgt_9_419, // sfix19_En18 
  input [18:0] Wgt_9_420, // sfix19_En18 
  input [18:0] Wgt_9_421, // sfix19_En18 
  input [18:0] Wgt_9_422, // sfix19_En18 
  input [18:0] Wgt_9_423, // sfix19_En18 
  input [18:0] Wgt_9_424, // sfix19_En18 
  input [18:0] Wgt_9_425, // sfix19_En18 
  input [18:0] Wgt_9_426, // sfix19_En18 
  input [18:0] Wgt_9_427, // sfix19_En18 
  input [18:0] Wgt_9_428, // sfix19_En18 
  input [18:0] Wgt_9_429, // sfix19_En18 
  input [18:0] Wgt_9_430, // sfix19_En18 
  input [18:0] Wgt_9_431, // sfix19_En18 
  input [18:0] Wgt_9_432, // sfix19_En18 
  input [18:0] Wgt_9_433, // sfix19_En18 
  input [18:0] Wgt_9_434, // sfix19_En18 
  input [18:0] Wgt_9_435, // sfix19_En18 
  input [18:0] Wgt_9_436, // sfix19_En18 
  input [18:0] Wgt_9_437, // sfix19_En18 
  input [18:0] Wgt_9_438, // sfix19_En18 
  input [18:0] Wgt_9_439, // sfix19_En18 
  input [18:0] Wgt_9_440, // sfix19_En18 
  input [18:0] Wgt_9_441, // sfix19_En18 
  input [18:0] Wgt_9_442, // sfix19_En18 
  input [18:0] Wgt_9_443, // sfix19_En18 
  input [18:0] Wgt_9_444, // sfix19_En18 
  input [18:0] Wgt_9_445, // sfix19_En18 
  input [18:0] Wgt_9_446, // sfix19_En18 
  input [18:0] Wgt_9_447, // sfix19_En18 
  input [18:0] Wgt_9_448, // sfix19_En18 
  input [18:0] Wgt_9_449, // sfix19_En18 
  input [18:0] Wgt_9_450, // sfix19_En18 
  input [18:0] Wgt_9_451, // sfix19_En18 
  input [18:0] Wgt_9_452, // sfix19_En18 
  input [18:0] Wgt_9_453, // sfix19_En18 
  input [18:0] Wgt_9_454, // sfix19_En18 
  input [18:0] Wgt_9_455, // sfix19_En18 
  input [18:0] Wgt_9_456, // sfix19_En18 
  input [18:0] Wgt_9_457, // sfix19_En18 
  input [18:0] Wgt_9_458, // sfix19_En18 
  input [18:0] Wgt_9_459, // sfix19_En18 
  input [18:0] Wgt_9_460, // sfix19_En18 
  input [18:0] Wgt_9_461, // sfix19_En18 
  input [18:0] Wgt_9_462, // sfix19_En18 
  input [18:0] Wgt_9_463, // sfix19_En18 
  input [18:0] Wgt_9_464, // sfix19_En18 
  input [18:0] Wgt_9_465, // sfix19_En18 
  input [18:0] Wgt_9_466, // sfix19_En18 
  input [18:0] Wgt_9_467, // sfix19_En18 
  input [18:0] Wgt_9_468, // sfix19_En18 
  input [18:0] Wgt_9_469, // sfix19_En18 
  input [18:0] Wgt_9_470, // sfix19_En18 
  input [18:0] Wgt_9_471, // sfix19_En18 
  input [18:0] Wgt_9_472, // sfix19_En18 
  input [18:0] Wgt_9_473, // sfix19_En18 
  input [18:0] Wgt_9_474, // sfix19_En18 
  input [18:0] Wgt_9_475, // sfix19_En18 
  input [18:0] Wgt_9_476, // sfix19_En18 
  input [18:0] Wgt_9_477, // sfix19_En18 
  input [18:0] Wgt_9_478, // sfix19_En18 
  input [18:0] Wgt_9_479, // sfix19_En18 
  input [18:0] Wgt_9_480, // sfix19_En18 
  input [18:0] Wgt_9_481, // sfix19_En18 
  input [18:0] Wgt_9_482, // sfix19_En18 
  input [18:0] Wgt_9_483, // sfix19_En18 
  input [18:0] Wgt_9_484, // sfix19_En18 
  input [18:0] Wgt_9_485, // sfix19_En18 
  input [18:0] Wgt_9_486, // sfix19_En18 
  input [18:0] Wgt_9_487, // sfix19_En18 
  input [18:0] Wgt_9_488, // sfix19_En18 
  input [18:0] Wgt_9_489, // sfix19_En18 
  input [18:0] Wgt_9_490, // sfix19_En18 
  input [18:0] Wgt_9_491, // sfix19_En18 
  input [18:0] Wgt_9_492, // sfix19_En18 
  input [18:0] Wgt_9_493, // sfix19_En18 
  input [18:0] Wgt_9_494, // sfix19_En18 
  input [18:0] Wgt_9_495, // sfix19_En18 
  input [18:0] Wgt_9_496, // sfix19_En18 
  input [18:0] Wgt_9_497, // sfix19_En18 
  input [18:0] Wgt_9_498, // sfix19_En18 
  input [18:0] Wgt_9_499, // sfix19_En18 
  input [18:0] Wgt_9_500, // sfix19_En18 
  input [18:0] Wgt_9_501, // sfix19_En18 
  input [18:0] Wgt_9_502, // sfix19_En18 
  input [18:0] Wgt_9_503, // sfix19_En18 
  input [18:0] Wgt_9_504, // sfix19_En18 
  input [18:0] Wgt_9_505, // sfix19_En18 
  input [18:0] Wgt_9_506, // sfix19_En18 
  input [18:0] Wgt_9_507, // sfix19_En18 
  input [18:0] Wgt_9_508, // sfix19_En18 
  input [18:0] Wgt_9_509, // sfix19_En18 
  input [18:0] Wgt_9_510, // sfix19_En18 
  input [18:0] Wgt_9_511, // sfix19_En18 
  input [18:0] Wgt_9_512, // sfix19_En18 
  input [18:0] Wgt_9_513, // sfix19_En18 
  input [18:0] Wgt_9_514, // sfix19_En18 
  input [18:0] Wgt_9_515, // sfix19_En18 
  input [18:0] Wgt_9_516, // sfix19_En18 
  input [18:0] Wgt_9_517, // sfix19_En18 
  input [18:0] Wgt_9_518, // sfix19_En18 
  input [18:0] Wgt_9_519, // sfix19_En18 
  input [18:0] Wgt_9_520, // sfix19_En18 
  input [18:0] Wgt_9_521, // sfix19_En18 
  input [18:0] Wgt_9_522, // sfix19_En18 
  input [18:0] Wgt_9_523, // sfix19_En18 
  input [18:0] Wgt_9_524, // sfix19_En18 
  input [18:0] Wgt_9_525, // sfix19_En18 
  input [18:0] Wgt_9_526, // sfix19_En18 
  input [18:0] Wgt_9_527, // sfix19_En18 
  input [18:0] Wgt_9_528, // sfix19_En18 
  input [18:0] Wgt_9_529, // sfix19_En18 
  input [18:0] Wgt_9_530, // sfix19_En18 
  input [18:0] Wgt_9_531, // sfix19_En18 
  input [18:0] Wgt_9_532, // sfix19_En18 
  input [18:0] Wgt_9_533, // sfix19_En18 
  input [18:0] Wgt_9_534, // sfix19_En18 
  input [18:0] Wgt_9_535, // sfix19_En18 
  input [18:0] Wgt_9_536, // sfix19_En18 
  input [18:0] Wgt_9_537, // sfix19_En18 
  input [18:0] Wgt_9_538, // sfix19_En18 
  input [18:0] Wgt_9_539, // sfix19_En18 
  input [18:0] Wgt_9_540, // sfix19_En18 
  input [18:0] Wgt_9_541, // sfix19_En18 
  input [18:0] Wgt_9_542, // sfix19_En18 
  input [18:0] Wgt_9_543, // sfix19_En18 
  input [18:0] Wgt_9_544, // sfix19_En18 
  input [18:0] Wgt_9_545, // sfix19_En18 
  input [18:0] Wgt_9_546, // sfix19_En18 
  input [18:0] Wgt_9_547, // sfix19_En18 
  input [18:0] Wgt_9_548, // sfix19_En18 
  input [18:0] Wgt_9_549, // sfix19_En18 
  input [18:0] Wgt_9_550, // sfix19_En18 
  input [18:0] Wgt_9_551, // sfix19_En18 
  input [18:0] Wgt_9_552, // sfix19_En18 
  input [18:0] Wgt_9_553, // sfix19_En18 
  input [18:0] Wgt_9_554, // sfix19_En18 
  input [18:0] Wgt_9_555, // sfix19_En18 
  input [18:0] Wgt_9_556, // sfix19_En18 
  input [18:0] Wgt_9_557, // sfix19_En18 
  input [18:0] Wgt_9_558, // sfix19_En18 
  input [18:0] Wgt_9_559, // sfix19_En18 
  input [18:0] Wgt_9_560, // sfix19_En18 
  input [18:0] Wgt_9_561, // sfix19_En18 
  input [18:0] Wgt_9_562, // sfix19_En18 
  input [18:0] Wgt_9_563, // sfix19_En18 
  input [18:0] Wgt_9_564, // sfix19_En18 
  input [18:0] Wgt_9_565, // sfix19_En18 
  input [18:0] Wgt_9_566, // sfix19_En18 
  input [18:0] Wgt_9_567, // sfix19_En18 
  input [18:0] Wgt_9_568, // sfix19_En18 
  input [18:0] Wgt_9_569, // sfix19_En18 
  input [18:0] Wgt_9_570, // sfix19_En18 
  input [18:0] Wgt_9_571, // sfix19_En18 
  input [18:0] Wgt_9_572, // sfix19_En18 
  input [18:0] Wgt_9_573, // sfix19_En18 
  input [18:0] Wgt_9_574, // sfix19_En18 
  input [18:0] Wgt_9_575, // sfix19_En18 
  input [18:0] Wgt_9_576, // sfix19_En18 
  input [18:0] Wgt_9_577, // sfix19_En18 
  input [18:0] Wgt_9_578, // sfix19_En18 
  input [18:0] Wgt_9_579, // sfix19_En18 
  input [18:0] Wgt_9_580, // sfix19_En18 
  input [18:0] Wgt_9_581, // sfix19_En18 
  input [18:0] Wgt_9_582, // sfix19_En18 
  input [18:0] Wgt_9_583, // sfix19_En18 
  input [18:0] Wgt_9_584, // sfix19_En18 
  input [18:0] Wgt_9_585, // sfix19_En18 
  input [18:0] Wgt_9_586, // sfix19_En18 
  input [18:0] Wgt_9_587, // sfix19_En18 
  input [18:0] Wgt_9_588, // sfix19_En18 
  input [18:0] Wgt_9_589, // sfix19_En18 
  input [18:0] Wgt_9_590, // sfix19_En18 
  input [18:0] Wgt_9_591, // sfix19_En18 
  input [18:0] Wgt_9_592, // sfix19_En18 
  input [18:0] Wgt_9_593, // sfix19_En18 
  input [18:0] Wgt_9_594, // sfix19_En18 
  input [18:0] Wgt_9_595, // sfix19_En18 
  input [18:0] Wgt_9_596, // sfix19_En18 
  input [18:0] Wgt_9_597, // sfix19_En18 
  input [18:0] Wgt_9_598, // sfix19_En18 
  input [18:0] Wgt_9_599, // sfix19_En18 
  input [18:0] Wgt_9_600, // sfix19_En18 
  input [18:0] Wgt_9_601, // sfix19_En18 
  input [18:0] Wgt_9_602, // sfix19_En18 
  input [18:0] Wgt_9_603, // sfix19_En18 
  input [18:0] Wgt_9_604, // sfix19_En18 
  input [18:0] Wgt_9_605, // sfix19_En18 
  input [18:0] Wgt_9_606, // sfix19_En18 
  input [18:0] Wgt_9_607, // sfix19_En18 
  input [18:0] Wgt_9_608, // sfix19_En18 
  input [18:0] Wgt_9_609, // sfix19_En18 
  input [18:0] Wgt_9_610, // sfix19_En18 
  input [18:0] Wgt_9_611, // sfix19_En18 
  input [18:0] Wgt_9_612, // sfix19_En18 
  input [18:0] Wgt_9_613, // sfix19_En18 
  input [18:0] Wgt_9_614, // sfix19_En18 
  input [18:0] Wgt_9_615, // sfix19_En18 
  input [18:0] Wgt_9_616, // sfix19_En18 
  input [18:0] Wgt_9_617, // sfix19_En18 
  input [18:0] Wgt_9_618, // sfix19_En18 
  input [18:0] Wgt_9_619, // sfix19_En18 
  input [18:0] Wgt_9_620, // sfix19_En18 
  input [18:0] Wgt_9_621, // sfix19_En18 
  input [18:0] Wgt_9_622, // sfix19_En18 
  input [18:0] Wgt_9_623, // sfix19_En18 
  input [18:0] Wgt_9_624, // sfix19_En18 
  input [18:0] Wgt_9_625, // sfix19_En18 
  input [18:0] Wgt_9_626, // sfix19_En18 
  input [18:0] Wgt_9_627, // sfix19_En18 
  input [18:0] Wgt_9_628, // sfix19_En18 
  input [18:0] Wgt_9_629, // sfix19_En18 
  input [18:0] Wgt_9_630, // sfix19_En18 
  input [18:0] Wgt_9_631, // sfix19_En18 
  input [18:0] Wgt_9_632, // sfix19_En18 
  input [18:0] Wgt_9_633, // sfix19_En18 
  input [18:0] Wgt_9_634, // sfix19_En18 
  input [18:0] Wgt_9_635, // sfix19_En18 
  input [18:0] Wgt_9_636, // sfix19_En18 
  input [18:0] Wgt_9_637, // sfix19_En18 
  input [18:0] Wgt_9_638, // sfix19_En18 
  input [18:0] Wgt_9_639, // sfix19_En18 
  input [18:0] Wgt_9_640, // sfix19_En18 
  input [18:0] Wgt_9_641, // sfix19_En18 
  input [18:0] Wgt_9_642, // sfix19_En18 
  input [18:0] Wgt_9_643, // sfix19_En18 
  input [18:0] Wgt_9_644, // sfix19_En18 
  input [18:0] Wgt_9_645, // sfix19_En18 
  input [18:0] Wgt_9_646, // sfix19_En18 
  input [18:0] Wgt_9_647, // sfix19_En18 
  input [18:0] Wgt_9_648, // sfix19_En18 
  input [18:0] Wgt_9_649, // sfix19_En18 
  input [18:0] Wgt_9_650, // sfix19_En18 
  input [18:0] Wgt_9_651, // sfix19_En18 
  input [18:0] Wgt_9_652, // sfix19_En18 
  input [18:0] Wgt_9_653, // sfix19_En18 
  input [18:0] Wgt_9_654, // sfix19_En18 
  input [18:0] Wgt_9_655, // sfix19_En18 
  input [18:0] Wgt_9_656, // sfix19_En18 
  input [18:0] Wgt_9_657, // sfix19_En18 
  input [18:0] Wgt_9_658, // sfix19_En18 
  input [18:0] Wgt_9_659, // sfix19_En18 
  input [18:0] Wgt_9_660, // sfix19_En18 
  input [18:0] Wgt_9_661, // sfix19_En18 
  input [18:0] Wgt_9_662, // sfix19_En18 
  input [18:0] Wgt_9_663, // sfix19_En18 
  input [18:0] Wgt_9_664, // sfix19_En18 
  input [18:0] Wgt_9_665, // sfix19_En18 
  input [18:0] Wgt_9_666, // sfix19_En18 
  input [18:0] Wgt_9_667, // sfix19_En18 
  input [18:0] Wgt_9_668, // sfix19_En18 
  input [18:0] Wgt_9_669, // sfix19_En18 
  input [18:0] Wgt_9_670, // sfix19_En18 
  input [18:0] Wgt_9_671, // sfix19_En18 
  input [18:0] Wgt_9_672, // sfix19_En18 
  input [18:0] Wgt_9_673, // sfix19_En18 
  input [18:0] Wgt_9_674, // sfix19_En18 
  input [18:0] Wgt_9_675, // sfix19_En18 
  input [18:0] Wgt_9_676, // sfix19_En18 
  input [18:0] Wgt_9_677, // sfix19_En18 
  input [18:0] Wgt_9_678, // sfix19_En18 
  input [18:0] Wgt_9_679, // sfix19_En18 
  input [18:0] Wgt_9_680, // sfix19_En18 
  input [18:0] Wgt_9_681, // sfix19_En18 
  input [18:0] Wgt_9_682, // sfix19_En18 
  input [18:0] Wgt_9_683, // sfix19_En18 
  input [18:0] Wgt_9_684, // sfix19_En18 
  input [18:0] Wgt_9_685, // sfix19_En18 
  input [18:0] Wgt_9_686, // sfix19_En18 
  input [18:0] Wgt_9_687, // sfix19_En18 
  input [18:0] Wgt_9_688, // sfix19_En18 
  input [18:0] Wgt_9_689, // sfix19_En18 
  input [18:0] Wgt_9_690, // sfix19_En18 
  input [18:0] Wgt_9_691, // sfix19_En18 
  input [18:0] Wgt_9_692, // sfix19_En18 
  input [18:0] Wgt_9_693, // sfix19_En18 
  input [18:0] Wgt_9_694, // sfix19_En18 
  input [18:0] Wgt_9_695, // sfix19_En18 
  input [18:0] Wgt_9_696, // sfix19_En18 
  input [18:0] Wgt_9_697, // sfix19_En18 
  input [18:0] Wgt_9_698, // sfix19_En18 
  input [18:0] Wgt_9_699, // sfix19_En18 
  input [18:0] Wgt_9_700, // sfix19_En18 
  input [18:0] Wgt_9_701, // sfix19_En18 
  input [18:0] Wgt_9_702, // sfix19_En18 
  input [18:0] Wgt_9_703, // sfix19_En18 
  input [18:0] Wgt_9_704, // sfix19_En18 
  input [18:0] Wgt_9_705, // sfix19_En18 
  input [18:0] Wgt_9_706, // sfix19_En18 
  input [18:0] Wgt_9_707, // sfix19_En18 
  input [18:0] Wgt_9_708, // sfix19_En18 
  input [18:0] Wgt_9_709, // sfix19_En18 
  input [18:0] Wgt_9_710, // sfix19_En18 
  input [18:0] Wgt_9_711, // sfix19_En18 
  input [18:0] Wgt_9_712, // sfix19_En18 
  input [18:0] Wgt_9_713, // sfix19_En18 
  input [18:0] Wgt_9_714, // sfix19_En18 
  input [18:0] Wgt_9_715, // sfix19_En18 
  input [18:0] Wgt_9_716, // sfix19_En18 
  input [18:0] Wgt_9_717, // sfix19_En18 
  input [18:0] Wgt_9_718, // sfix19_En18 
  input [18:0] Wgt_9_719, // sfix19_En18 
  input [18:0] Wgt_9_720, // sfix19_En18 
  input [18:0] Wgt_9_721, // sfix19_En18 
  input [18:0] Wgt_9_722, // sfix19_En18 
  input [18:0] Wgt_9_723, // sfix19_En18 
  input [18:0] Wgt_9_724, // sfix19_En18 
  input [18:0] Wgt_9_725, // sfix19_En18 
  input [18:0] Wgt_9_726, // sfix19_En18 
  input [18:0] Wgt_9_727, // sfix19_En18 
  input [18:0] Wgt_9_728, // sfix19_En18 
  input [18:0] Wgt_9_729, // sfix19_En18 
  input [18:0] Wgt_9_730, // sfix19_En18 
  input [18:0] Wgt_9_731, // sfix19_En18 
  input [18:0] Wgt_9_732, // sfix19_En18 
  input [18:0] Wgt_9_733, // sfix19_En18 
  input [18:0] Wgt_9_734, // sfix19_En18 
  input [18:0] Wgt_9_735, // sfix19_En18 
  input [18:0] Wgt_9_736, // sfix19_En18 
  input [18:0] Wgt_9_737, // sfix19_En18 
  input [18:0] Wgt_9_738, // sfix19_En18 
  input [18:0] Wgt_9_739, // sfix19_En18 
  input [18:0] Wgt_9_740, // sfix19_En18 
  input [18:0] Wgt_9_741, // sfix19_En18 
  input [18:0] Wgt_9_742, // sfix19_En18 
  input [18:0] Wgt_9_743, // sfix19_En18 
  input [18:0] Wgt_9_744, // sfix19_En18 
  input [18:0] Wgt_9_745, // sfix19_En18 
  input [18:0] Wgt_9_746, // sfix19_En18 
  input [18:0] Wgt_9_747, // sfix19_En18 
  input [18:0] Wgt_9_748, // sfix19_En18 
  input [18:0] Wgt_9_749, // sfix19_En18 
  input [18:0] Wgt_9_750, // sfix19_En18 
  input [18:0] Wgt_9_751, // sfix19_En18 
  input [18:0] Wgt_9_752, // sfix19_En18 
  input [18:0] Wgt_9_753, // sfix19_En18 
  input [18:0] Wgt_9_754, // sfix19_En18 
  input [18:0] Wgt_9_755, // sfix19_En18 
  input [18:0] Wgt_9_756, // sfix19_En18 
  input [18:0] Wgt_9_757, // sfix19_En18 
  input [18:0] Wgt_9_758, // sfix19_En18 
  input [18:0] Wgt_9_759, // sfix19_En18 
  input [18:0] Wgt_9_760, // sfix19_En18 
  input [18:0] Wgt_9_761, // sfix19_En18 
  input [18:0] Wgt_9_762, // sfix19_En18 
  input [18:0] Wgt_9_763, // sfix19_En18 
  input [18:0] Wgt_9_764, // sfix19_En18 
  input [18:0] Wgt_9_765, // sfix19_En18 
  input [18:0] Wgt_9_766, // sfix19_En18 
  input [18:0] Wgt_9_767, // sfix19_En18 
  input [18:0] Wgt_9_768, // sfix19_En18 
  input [18:0] Wgt_9_769, // sfix19_En18 
  input [18:0] Wgt_9_770, // sfix19_En18 
  input [18:0] Wgt_9_771, // sfix19_En18 
  input [18:0] Wgt_9_772, // sfix19_En18 
  input [18:0] Wgt_9_773, // sfix19_En18 
  input [18:0] Wgt_9_774, // sfix19_En18 
  input [18:0] Wgt_9_775, // sfix19_En18 
  input [18:0] Wgt_9_776, // sfix19_En18 
  input [18:0] Wgt_9_777, // sfix19_En18 
  input [18:0] Wgt_9_778, // sfix19_En18 
  input [18:0] Wgt_9_779, // sfix19_En18 
  input [18:0] Wgt_9_780, // sfix19_En18 
  input [18:0] Wgt_9_781, // sfix19_En18 
  input [18:0] Wgt_9_782, // sfix19_En18 
  input [18:0] Wgt_9_783, // sfix19_En18 
  input [18:0] Wgt_9_784, // sfix19_En18 
  input [9:0] Pix_0, // sfix10_En0 
 input [9:0] Pix_1, // sfix10_En0 
    input [9:0] Pix_2, // sfix10_En0 
    input [9:0] Pix_3, // sfix10_En0 
    input [9:0] Pix_4, // sfix10_En0 
    input [9:0] Pix_5, // sfix10_En0 
    input [9:0] Pix_6, // sfix10_En0 
    input [9:0] Pix_7, // sfix10_En0 
    input [9:0] Pix_8, // sfix10_En0 
    input [9:0] Pix_9, // sfix10_En0 
    input [9:0] Pix_10, // sfix10_En0 
    input [9:0] Pix_11, // sfix10_En0 
    input [9:0] Pix_12, // sfix10_En0 
    input [9:0] Pix_13, // sfix10_En0 
    input [9:0] Pix_14, // sfix10_En0 
    input [9:0] Pix_15, // sfix10_En0 
    input [9:0] Pix_16, // sfix10_En0 
    input [9:0] Pix_17, // sfix10_En0 
    input [9:0] Pix_18, // sfix10_En0 
    input [9:0] Pix_19, // sfix10_En0 
    input [9:0] Pix_20, // sfix10_En0 
    input [9:0] Pix_21, // sfix10_En0 
    input [9:0] Pix_22, // sfix10_En0 
    input [9:0] Pix_23, // sfix10_En0 
    input [9:0] Pix_24, // sfix10_En0 
    input [9:0] Pix_25, // sfix10_En0 
    input [9:0] Pix_26, // sfix10_En0 
    input [9:0] Pix_27, // sfix10_En0 
    input [9:0] Pix_28, // sfix10_En0 
    input [9:0] Pix_29, // sfix10_En0 
    input [9:0] Pix_30, // sfix10_En0 
    input [9:0] Pix_31, // sfix10_En0 
    input [9:0] Pix_32, // sfix10_En0 
    input [9:0] Pix_33, // sfix10_En0 
    input [9:0] Pix_34, // sfix10_En0 
    input [9:0] Pix_35, // sfix10_En0 
    input [9:0] Pix_36, // sfix10_En0 
    input [9:0] Pix_37, // sfix10_En0 
    input [9:0] Pix_38, // sfix10_En0 
    input [9:0] Pix_39, // sfix10_En0 
    input [9:0] Pix_40, // sfix10_En0 
    input [9:0] Pix_41, // sfix10_En0 
    input [9:0] Pix_42, // sfix10_En0 
    input [9:0] Pix_43, // sfix10_En0 
    input [9:0] Pix_44, // sfix10_En0 
    input [9:0] Pix_45, // sfix10_En0 
    input [9:0] Pix_46, // sfix10_En0 
    input [9:0] Pix_47, // sfix10_En0 
    input [9:0] Pix_48, // sfix10_En0 
    input [9:0] Pix_49, // sfix10_En0 
    input [9:0] Pix_50, // sfix10_En0 
    input [9:0] Pix_51, // sfix10_En0 
    input [9:0] Pix_52, // sfix10_En0 
    input [9:0] Pix_53, // sfix10_En0 
    input [9:0] Pix_54, // sfix10_En0 
    input [9:0] Pix_55, // sfix10_En0 
    input [9:0] Pix_56, // sfix10_En0 
    input [9:0] Pix_57, // sfix10_En0 
    input [9:0] Pix_58, // sfix10_En0 
    input [9:0] Pix_59, // sfix10_En0 
    input [9:0] Pix_60, // sfix10_En0 
    input [9:0] Pix_61, // sfix10_En0 
    input [9:0] Pix_62, // sfix10_En0 
    input [9:0] Pix_63, // sfix10_En0 
    input [9:0] Pix_64, // sfix10_En0 
    input [9:0] Pix_65, // sfix10_En0 
    input [9:0] Pix_66, // sfix10_En0 
    input [9:0] Pix_67, // sfix10_En0 
    input [9:0] Pix_68, // sfix10_En0 
    input [9:0] Pix_69, // sfix10_En0 
    input [9:0] Pix_70, // sfix10_En0 
    input [9:0] Pix_71, // sfix10_En0 
    input [9:0] Pix_72, // sfix10_En0 
    input [9:0] Pix_73, // sfix10_En0 
    input [9:0] Pix_74, // sfix10_En0 
    input [9:0] Pix_75, // sfix10_En0 
    input [9:0] Pix_76, // sfix10_En0 
    input [9:0] Pix_77, // sfix10_En0 
    input [9:0] Pix_78, // sfix10_En0 
    input [9:0] Pix_79, // sfix10_En0 
    input [9:0] Pix_80, // sfix10_En0 
    input [9:0] Pix_81, // sfix10_En0 
    input [9:0] Pix_82, // sfix10_En0 
    input [9:0] Pix_83, // sfix10_En0 
    input [9:0] Pix_84, // sfix10_En0 
    input [9:0] Pix_85, // sfix10_En0 
    input [9:0] Pix_86, // sfix10_En0 
    input [9:0] Pix_87, // sfix10_En0 
    input [9:0] Pix_88, // sfix10_En0 
    input [9:0] Pix_89, // sfix10_En0 
    input [9:0] Pix_90, // sfix10_En0 
    input [9:0] Pix_91, // sfix10_En0 
    input [9:0] Pix_92, // sfix10_En0 
    input [9:0] Pix_93, // sfix10_En0 
    input [9:0] Pix_94, // sfix10_En0 
    input [9:0] Pix_95, // sfix10_En0 
    input [9:0] Pix_96, // sfix10_En0 
    input [9:0] Pix_97, // sfix10_En0 
    input [9:0] Pix_98, // sfix10_En0 
    input [9:0] Pix_99, // sfix10_En0 
    input [9:0] Pix_100, // sfix10_En0 
    input [9:0] Pix_101, // sfix10_En0 
    input [9:0] Pix_102, // sfix10_En0 
    input [9:0] Pix_103, // sfix10_En0 
    input [9:0] Pix_104, // sfix10_En0 
    input [9:0] Pix_105, // sfix10_En0 
    input [9:0] Pix_106, // sfix10_En0 
    input [9:0] Pix_107, // sfix10_En0 
    input [9:0] Pix_108, // sfix10_En0 
    input [9:0] Pix_109, // sfix10_En0 
    input [9:0] Pix_110, // sfix10_En0 
    input [9:0] Pix_111, // sfix10_En0 
    input [9:0] Pix_112, // sfix10_En0 
    input [9:0] Pix_113, // sfix10_En0 
    input [9:0] Pix_114, // sfix10_En0 
    input [9:0] Pix_115, // sfix10_En0 
    input [9:0] Pix_116, // sfix10_En0 
    input [9:0] Pix_117, // sfix10_En0 
    input [9:0] Pix_118, // sfix10_En0 
    input [9:0] Pix_119, // sfix10_En0 
    input [9:0] Pix_120, // sfix10_En0 
    input [9:0] Pix_121, // sfix10_En0 
    input [9:0] Pix_122, // sfix10_En0 
    input [9:0] Pix_123, // sfix10_En0 
    input [9:0] Pix_124, // sfix10_En0 
    input [9:0] Pix_125, // sfix10_En0 
    input [9:0] Pix_126, // sfix10_En0 
    input [9:0] Pix_127, // sfix10_En0 
    input [9:0] Pix_128, // sfix10_En0 
    input [9:0] Pix_129, // sfix10_En0 
    input [9:0] Pix_130, // sfix10_En0 
    input [9:0] Pix_131, // sfix10_En0 
    input [9:0] Pix_132, // sfix10_En0 
    input [9:0] Pix_133, // sfix10_En0 
    input [9:0] Pix_134, // sfix10_En0 
    input [9:0] Pix_135, // sfix10_En0 
    input [9:0] Pix_136, // sfix10_En0 
    input [9:0] Pix_137, // sfix10_En0 
    input [9:0] Pix_138, // sfix10_En0 
    input [9:0] Pix_139, // sfix10_En0 
    input [9:0] Pix_140, // sfix10_En0 
    input [9:0] Pix_141, // sfix10_En0 
    input [9:0] Pix_142, // sfix10_En0 
    input [9:0] Pix_143, // sfix10_En0 
    input [9:0] Pix_144, // sfix10_En0 
    input [9:0] Pix_145, // sfix10_En0 
    input [9:0] Pix_146, // sfix10_En0 
    input [9:0] Pix_147, // sfix10_En0 
    input [9:0] Pix_148, // sfix10_En0 
    input [9:0] Pix_149, // sfix10_En0 
    input [9:0] Pix_150, // sfix10_En0 
    input [9:0] Pix_151, // sfix10_En0 
    input [9:0] Pix_152, // sfix10_En0 
    input [9:0] Pix_153, // sfix10_En0 
    input [9:0] Pix_154, // sfix10_En0 
    input [9:0] Pix_155, // sfix10_En0 
    input [9:0] Pix_156, // sfix10_En0 
    input [9:0] Pix_157, // sfix10_En0 
    input [9:0] Pix_158, // sfix10_En0 
    input [9:0] Pix_159, // sfix10_En0 
    input [9:0] Pix_160, // sfix10_En0 
    input [9:0] Pix_161, // sfix10_En0 
    input [9:0] Pix_162, // sfix10_En0 
    input [9:0] Pix_163, // sfix10_En0 
    input [9:0] Pix_164, // sfix10_En0 
    input [9:0] Pix_165, // sfix10_En0 
    input [9:0] Pix_166, // sfix10_En0 
    input [9:0] Pix_167, // sfix10_En0 
    input [9:0] Pix_168, // sfix10_En0 
    input [9:0] Pix_169, // sfix10_En0 
    input [9:0] Pix_170, // sfix10_En0 
    input [9:0] Pix_171, // sfix10_En0 
    input [9:0] Pix_172, // sfix10_En0 
    input [9:0] Pix_173, // sfix10_En0 
    input [9:0] Pix_174, // sfix10_En0 
    input [9:0] Pix_175, // sfix10_En0 
    input [9:0] Pix_176, // sfix10_En0 
    input [9:0] Pix_177, // sfix10_En0 
    input [9:0] Pix_178, // sfix10_En0 
    input [9:0] Pix_179, // sfix10_En0 
    input [9:0] Pix_180, // sfix10_En0 
    input [9:0] Pix_181, // sfix10_En0 
    input [9:0] Pix_182, // sfix10_En0 
    input [9:0] Pix_183, // sfix10_En0 
    input [9:0] Pix_184, // sfix10_En0 
    input [9:0] Pix_185, // sfix10_En0 
    input [9:0] Pix_186, // sfix10_En0 
    input [9:0] Pix_187, // sfix10_En0 
    input [9:0] Pix_188, // sfix10_En0 
    input [9:0] Pix_189, // sfix10_En0 
    input [9:0] Pix_190, // sfix10_En0 
    input [9:0] Pix_191, // sfix10_En0 
    input [9:0] Pix_192, // sfix10_En0 
    input [9:0] Pix_193, // sfix10_En0 
    input [9:0] Pix_194, // sfix10_En0 
    input [9:0] Pix_195, // sfix10_En0 
    input [9:0] Pix_196, // sfix10_En0 
    input [9:0] Pix_197, // sfix10_En0 
    input [9:0] Pix_198, // sfix10_En0 
    input [9:0] Pix_199, // sfix10_En0 
    input [9:0] Pix_200, // sfix10_En0 
    input [9:0] Pix_201, // sfix10_En0 
    input [9:0] Pix_202, // sfix10_En0 
    input [9:0] Pix_203, // sfix10_En0 
    input [9:0] Pix_204, // sfix10_En0 
    input [9:0] Pix_205, // sfix10_En0 
    input [9:0] Pix_206, // sfix10_En0 
    input [9:0] Pix_207, // sfix10_En0 
    input [9:0] Pix_208, // sfix10_En0 
    input [9:0] Pix_209, // sfix10_En0 
    input [9:0] Pix_210, // sfix10_En0 
    input [9:0] Pix_211, // sfix10_En0 
    input [9:0] Pix_212, // sfix10_En0 
    input [9:0] Pix_213, // sfix10_En0 
    input [9:0] Pix_214, // sfix10_En0 
    input [9:0] Pix_215, // sfix10_En0 
    input [9:0] Pix_216, // sfix10_En0 
    input [9:0] Pix_217, // sfix10_En0 
    input [9:0] Pix_218, // sfix10_En0 
    input [9:0] Pix_219, // sfix10_En0 
    input [9:0] Pix_220, // sfix10_En0 
    input [9:0] Pix_221, // sfix10_En0 
    input [9:0] Pix_222, // sfix10_En0 
    input [9:0] Pix_223, // sfix10_En0 
    input [9:0] Pix_224, // sfix10_En0 
    input [9:0] Pix_225, // sfix10_En0 
    input [9:0] Pix_226, // sfix10_En0 
    input [9:0] Pix_227, // sfix10_En0 
    input [9:0] Pix_228, // sfix10_En0 
    input [9:0] Pix_229, // sfix10_En0 
    input [9:0] Pix_230, // sfix10_En0 
    input [9:0] Pix_231, // sfix10_En0 
    input [9:0] Pix_232, // sfix10_En0 
    input [9:0] Pix_233, // sfix10_En0 
    input [9:0] Pix_234, // sfix10_En0 
    input [9:0] Pix_235, // sfix10_En0 
    input [9:0] Pix_236, // sfix10_En0 
    input [9:0] Pix_237, // sfix10_En0 
    input [9:0] Pix_238, // sfix10_En0 
    input [9:0] Pix_239, // sfix10_En0 
    input [9:0] Pix_240, // sfix10_En0 
    input [9:0] Pix_241, // sfix10_En0 
    input [9:0] Pix_242, // sfix10_En0 
    input [9:0] Pix_243, // sfix10_En0 
    input [9:0] Pix_244, // sfix10_En0 
    input [9:0] Pix_245, // sfix10_En0 
    input [9:0] Pix_246, // sfix10_En0 
    input [9:0] Pix_247, // sfix10_En0 
    input [9:0] Pix_248, // sfix10_En0 
    input [9:0] Pix_249, // sfix10_En0 
    input [9:0] Pix_250, // sfix10_En0 
    input [9:0] Pix_251, // sfix10_En0 
    input [9:0] Pix_252, // sfix10_En0 
    input [9:0] Pix_253, // sfix10_En0 
    input [9:0] Pix_254, // sfix10_En0 
    input [9:0] Pix_255, // sfix10_En0 
    input [9:0] Pix_256, // sfix10_En0 
    input [9:0] Pix_257, // sfix10_En0 
    input [9:0] Pix_258, // sfix10_En0 
    input [9:0] Pix_259, // sfix10_En0 
    input [9:0] Pix_260, // sfix10_En0 
    input [9:0] Pix_261, // sfix10_En0 
    input [9:0] Pix_262, // sfix10_En0 
    input [9:0] Pix_263, // sfix10_En0 
    input [9:0] Pix_264, // sfix10_En0 
    input [9:0] Pix_265, // sfix10_En0 
    input [9:0] Pix_266, // sfix10_En0 
    input [9:0] Pix_267, // sfix10_En0 
    input [9:0] Pix_268, // sfix10_En0 
    input [9:0] Pix_269, // sfix10_En0 
    input [9:0] Pix_270, // sfix10_En0 
    input [9:0] Pix_271, // sfix10_En0 
    input [9:0] Pix_272, // sfix10_En0 
    input [9:0] Pix_273, // sfix10_En0 
    input [9:0] Pix_274, // sfix10_En0 
    input [9:0] Pix_275, // sfix10_En0 
    input [9:0] Pix_276, // sfix10_En0 
    input [9:0] Pix_277, // sfix10_En0 
    input [9:0] Pix_278, // sfix10_En0 
    input [9:0] Pix_279, // sfix10_En0 
    input [9:0] Pix_280, // sfix10_En0 
    input [9:0] Pix_281, // sfix10_En0 
    input [9:0] Pix_282, // sfix10_En0 
    input [9:0] Pix_283, // sfix10_En0 
    input [9:0] Pix_284, // sfix10_En0 
    input [9:0] Pix_285, // sfix10_En0 
    input [9:0] Pix_286, // sfix10_En0 
    input [9:0] Pix_287, // sfix10_En0 
    input [9:0] Pix_288, // sfix10_En0 
    input [9:0] Pix_289, // sfix10_En0 
    input [9:0] Pix_290, // sfix10_En0 
    input [9:0] Pix_291, // sfix10_En0 
    input [9:0] Pix_292, // sfix10_En0 
    input [9:0] Pix_293, // sfix10_En0 
    input [9:0] Pix_294, // sfix10_En0 
    input [9:0] Pix_295, // sfix10_En0 
    input [9:0] Pix_296, // sfix10_En0 
    input [9:0] Pix_297, // sfix10_En0 
    input [9:0] Pix_298, // sfix10_En0 
    input [9:0] Pix_299, // sfix10_En0 
    input [9:0] Pix_300, // sfix10_En0 
    input [9:0] Pix_301, // sfix10_En0 
    input [9:0] Pix_302, // sfix10_En0 
    input [9:0] Pix_303, // sfix10_En0 
    input [9:0] Pix_304, // sfix10_En0 
    input [9:0] Pix_305, // sfix10_En0 
    input [9:0] Pix_306, // sfix10_En0 
    input [9:0] Pix_307, // sfix10_En0 
    input [9:0] Pix_308, // sfix10_En0 
    input [9:0] Pix_309, // sfix10_En0 
    input [9:0] Pix_310, // sfix10_En0 
    input [9:0] Pix_311, // sfix10_En0 
    input [9:0] Pix_312, // sfix10_En0 
    input [9:0] Pix_313, // sfix10_En0 
    input [9:0] Pix_314, // sfix10_En0 
    input [9:0] Pix_315, // sfix10_En0 
    input [9:0] Pix_316, // sfix10_En0 
    input [9:0] Pix_317, // sfix10_En0 
    input [9:0] Pix_318, // sfix10_En0 
    input [9:0] Pix_319, // sfix10_En0 
    input [9:0] Pix_320, // sfix10_En0 
    input [9:0] Pix_321, // sfix10_En0 
    input [9:0] Pix_322, // sfix10_En0 
    input [9:0] Pix_323, // sfix10_En0 
    input [9:0] Pix_324, // sfix10_En0 
    input [9:0] Pix_325, // sfix10_En0 
    input [9:0] Pix_326, // sfix10_En0 
    input [9:0] Pix_327, // sfix10_En0 
    input [9:0] Pix_328, // sfix10_En0 
    input [9:0] Pix_329, // sfix10_En0 
    input [9:0] Pix_330, // sfix10_En0 
    input [9:0] Pix_331, // sfix10_En0 
    input [9:0] Pix_332, // sfix10_En0 
    input [9:0] Pix_333, // sfix10_En0 
    input [9:0] Pix_334, // sfix10_En0 
    input [9:0] Pix_335, // sfix10_En0 
    input [9:0] Pix_336, // sfix10_En0 
    input [9:0] Pix_337, // sfix10_En0 
    input [9:0] Pix_338, // sfix10_En0 
    input [9:0] Pix_339, // sfix10_En0 
    input [9:0] Pix_340, // sfix10_En0 
    input [9:0] Pix_341, // sfix10_En0 
    input [9:0] Pix_342, // sfix10_En0 
    input [9:0] Pix_343, // sfix10_En0 
    input [9:0] Pix_344, // sfix10_En0 
    input [9:0] Pix_345, // sfix10_En0 
    input [9:0] Pix_346, // sfix10_En0 
    input [9:0] Pix_347, // sfix10_En0 
    input [9:0] Pix_348, // sfix10_En0 
    input [9:0] Pix_349, // sfix10_En0 
    input [9:0] Pix_350, // sfix10_En0 
    input [9:0] Pix_351, // sfix10_En0 
    input [9:0] Pix_352, // sfix10_En0 
    input [9:0] Pix_353, // sfix10_En0 
    input [9:0] Pix_354, // sfix10_En0 
    input [9:0] Pix_355, // sfix10_En0 
    input [9:0] Pix_356, // sfix10_En0 
    input [9:0] Pix_357, // sfix10_En0 
    input [9:0] Pix_358, // sfix10_En0 
    input [9:0] Pix_359, // sfix10_En0 
    input [9:0] Pix_360, // sfix10_En0 
    input [9:0] Pix_361, // sfix10_En0 
    input [9:0] Pix_362, // sfix10_En0 
    input [9:0] Pix_363, // sfix10_En0 
    input [9:0] Pix_364, // sfix10_En0 
    input [9:0] Pix_365, // sfix10_En0 
    input [9:0] Pix_366, // sfix10_En0 
    input [9:0] Pix_367, // sfix10_En0 
    input [9:0] Pix_368, // sfix10_En0 
    input [9:0] Pix_369, // sfix10_En0 
    input [9:0] Pix_370, // sfix10_En0 
    input [9:0] Pix_371, // sfix10_En0 
    input [9:0] Pix_372, // sfix10_En0 
    input [9:0] Pix_373, // sfix10_En0 
    input [9:0] Pix_374, // sfix10_En0 
    input [9:0] Pix_375, // sfix10_En0 
    input [9:0] Pix_376, // sfix10_En0 
    input [9:0] Pix_377, // sfix10_En0 
    input [9:0] Pix_378, // sfix10_En0 
    input [9:0] Pix_379, // sfix10_En0 
    input [9:0] Pix_380, // sfix10_En0 
    input [9:0] Pix_381, // sfix10_En0 
    input [9:0] Pix_382, // sfix10_En0 
    input [9:0] Pix_383, // sfix10_En0 
    input [9:0] Pix_384, // sfix10_En0 
    input [9:0] Pix_385, // sfix10_En0 
    input [9:0] Pix_386, // sfix10_En0 
    input [9:0] Pix_387, // sfix10_En0 
    input [9:0] Pix_388, // sfix10_En0 
    input [9:0] Pix_389, // sfix10_En0 
    input [9:0] Pix_390, // sfix10_En0 
    input [9:0] Pix_391, // sfix10_En0 
    input [9:0] Pix_392, // sfix10_En0 
    input [9:0] Pix_393, // sfix10_En0 
    input [9:0] Pix_394, // sfix10_En0 
    input [9:0] Pix_395, // sfix10_En0 
    input [9:0] Pix_396, // sfix10_En0 
    input [9:0] Pix_397, // sfix10_En0 
    input [9:0] Pix_398, // sfix10_En0 
    input [9:0] Pix_399, // sfix10_En0 
    input [9:0] Pix_400, // sfix10_En0 
    input [9:0] Pix_401, // sfix10_En0 
    input [9:0] Pix_402, // sfix10_En0 
    input [9:0] Pix_403, // sfix10_En0 
    input [9:0] Pix_404, // sfix10_En0 
    input [9:0] Pix_405, // sfix10_En0 
    input [9:0] Pix_406, // sfix10_En0 
    input [9:0] Pix_407, // sfix10_En0 
    input [9:0] Pix_408, // sfix10_En0 
    input [9:0] Pix_409, // sfix10_En0 
    input [9:0] Pix_410, // sfix10_En0 
    input [9:0] Pix_411, // sfix10_En0 
    input [9:0] Pix_412, // sfix10_En0 
    input [9:0] Pix_413, // sfix10_En0 
    input [9:0] Pix_414, // sfix10_En0 
    input [9:0] Pix_415, // sfix10_En0 
    input [9:0] Pix_416, // sfix10_En0 
    input [9:0] Pix_417, // sfix10_En0 
    input [9:0] Pix_418, // sfix10_En0 
    input [9:0] Pix_419, // sfix10_En0 
    input [9:0] Pix_420, // sfix10_En0 
    input [9:0] Pix_421, // sfix10_En0 
    input [9:0] Pix_422, // sfix10_En0 
    input [9:0] Pix_423, // sfix10_En0 
    input [9:0] Pix_424, // sfix10_En0 
    input [9:0] Pix_425, // sfix10_En0 
    input [9:0] Pix_426, // sfix10_En0 
    input [9:0] Pix_427, // sfix10_En0 
    input [9:0] Pix_428, // sfix10_En0 
    input [9:0] Pix_429, // sfix10_En0 
    input [9:0] Pix_430, // sfix10_En0 
    input [9:0] Pix_431, // sfix10_En0 
    input [9:0] Pix_432, // sfix10_En0 
    input [9:0] Pix_433, // sfix10_En0 
    input [9:0] Pix_434, // sfix10_En0 
    input [9:0] Pix_435, // sfix10_En0 
    input [9:0] Pix_436, // sfix10_En0 
    input [9:0] Pix_437, // sfix10_En0 
    input [9:0] Pix_438, // sfix10_En0 
    input [9:0] Pix_439, // sfix10_En0 
    input [9:0] Pix_440, // sfix10_En0 
    input [9:0] Pix_441, // sfix10_En0 
    input [9:0] Pix_442, // sfix10_En0 
    input [9:0] Pix_443, // sfix10_En0 
    input [9:0] Pix_444, // sfix10_En0 
    input [9:0] Pix_445, // sfix10_En0 
    input [9:0] Pix_446, // sfix10_En0 
    input [9:0] Pix_447, // sfix10_En0 
    input [9:0] Pix_448, // sfix10_En0 
    input [9:0] Pix_449, // sfix10_En0 
    input [9:0] Pix_450, // sfix10_En0 
    input [9:0] Pix_451, // sfix10_En0 
    input [9:0] Pix_452, // sfix10_En0 
    input [9:0] Pix_453, // sfix10_En0 
    input [9:0] Pix_454, // sfix10_En0 
    input [9:0] Pix_455, // sfix10_En0 
    input [9:0] Pix_456, // sfix10_En0 
    input [9:0] Pix_457, // sfix10_En0 
    input [9:0] Pix_458, // sfix10_En0 
    input [9:0] Pix_459, // sfix10_En0 
    input [9:0] Pix_460, // sfix10_En0 
    input [9:0] Pix_461, // sfix10_En0 
    input [9:0] Pix_462, // sfix10_En0 
    input [9:0] Pix_463, // sfix10_En0 
    input [9:0] Pix_464, // sfix10_En0 
    input [9:0] Pix_465, // sfix10_En0 
    input [9:0] Pix_466, // sfix10_En0 
    input [9:0] Pix_467, // sfix10_En0 
    input [9:0] Pix_468, // sfix10_En0 
    input [9:0] Pix_469, // sfix10_En0 
    input [9:0] Pix_470, // sfix10_En0 
    input [9:0] Pix_471, // sfix10_En0 
    input [9:0] Pix_472, // sfix10_En0 
    input [9:0] Pix_473, // sfix10_En0 
    input [9:0] Pix_474, // sfix10_En0 
    input [9:0] Pix_475, // sfix10_En0 
    input [9:0] Pix_476, // sfix10_En0 
    input [9:0] Pix_477, // sfix10_En0 
    input [9:0] Pix_478, // sfix10_En0 
    input [9:0] Pix_479, // sfix10_En0 
    input [9:0] Pix_480, // sfix10_En0 
    input [9:0] Pix_481, // sfix10_En0 
    input [9:0] Pix_482, // sfix10_En0 
    input [9:0] Pix_483, // sfix10_En0 
    input [9:0] Pix_484, // sfix10_En0 
    input [9:0] Pix_485, // sfix10_En0 
    input [9:0] Pix_486, // sfix10_En0 
    input [9:0] Pix_487, // sfix10_En0 
    input [9:0] Pix_488, // sfix10_En0 
    input [9:0] Pix_489, // sfix10_En0 
    input [9:0] Pix_490, // sfix10_En0 
    input [9:0] Pix_491, // sfix10_En0 
    input [9:0] Pix_492, // sfix10_En0 
    input [9:0] Pix_493, // sfix10_En0 
    input [9:0] Pix_494, // sfix10_En0 
    input [9:0] Pix_495, // sfix10_En0 
    input [9:0] Pix_496, // sfix10_En0 
    input [9:0] Pix_497, // sfix10_En0 
    input [9:0] Pix_498, // sfix10_En0 
    input [9:0] Pix_499, // sfix10_En0 
    input [9:0] Pix_500, // sfix10_En0 
    input [9:0] Pix_501, // sfix10_En0 
    input [9:0] Pix_502, // sfix10_En0 
    input [9:0] Pix_503, // sfix10_En0 
    input [9:0] Pix_504, // sfix10_En0 
    input [9:0] Pix_505, // sfix10_En0 
    input [9:0] Pix_506, // sfix10_En0 
    input [9:0] Pix_507, // sfix10_En0 
    input [9:0] Pix_508, // sfix10_En0 
    input [9:0] Pix_509, // sfix10_En0 
    input [9:0] Pix_510, // sfix10_En0 
    input [9:0] Pix_511, // sfix10_En0 
    input [9:0] Pix_512, // sfix10_En0 
    input [9:0] Pix_513, // sfix10_En0 
    input [9:0] Pix_514, // sfix10_En0 
    input [9:0] Pix_515, // sfix10_En0 
    input [9:0] Pix_516, // sfix10_En0 
    input [9:0] Pix_517, // sfix10_En0 
    input [9:0] Pix_518, // sfix10_En0 
    input [9:0] Pix_519, // sfix10_En0 
    input [9:0] Pix_520, // sfix10_En0 
    input [9:0] Pix_521, // sfix10_En0 
    input [9:0] Pix_522, // sfix10_En0 
    input [9:0] Pix_523, // sfix10_En0 
    input [9:0] Pix_524, // sfix10_En0 
    input [9:0] Pix_525, // sfix10_En0 
    input [9:0] Pix_526, // sfix10_En0 
    input [9:0] Pix_527, // sfix10_En0 
    input [9:0] Pix_528, // sfix10_En0 
    input [9:0] Pix_529, // sfix10_En0 
    input [9:0] Pix_530, // sfix10_En0 
    input [9:0] Pix_531, // sfix10_En0 
    input [9:0] Pix_532, // sfix10_En0 
    input [9:0] Pix_533, // sfix10_En0 
    input [9:0] Pix_534, // sfix10_En0 
    input [9:0] Pix_535, // sfix10_En0 
    input [9:0] Pix_536, // sfix10_En0 
    input [9:0] Pix_537, // sfix10_En0 
    input [9:0] Pix_538, // sfix10_En0 
    input [9:0] Pix_539, // sfix10_En0 
    input [9:0] Pix_540, // sfix10_En0 
    input [9:0] Pix_541, // sfix10_En0 
    input [9:0] Pix_542, // sfix10_En0 
    input [9:0] Pix_543, // sfix10_En0 
    input [9:0] Pix_544, // sfix10_En0 
    input [9:0] Pix_545, // sfix10_En0 
    input [9:0] Pix_546, // sfix10_En0 
    input [9:0] Pix_547, // sfix10_En0 
    input [9:0] Pix_548, // sfix10_En0 
    input [9:0] Pix_549, // sfix10_En0 
    input [9:0] Pix_550, // sfix10_En0 
    input [9:0] Pix_551, // sfix10_En0 
    input [9:0] Pix_552, // sfix10_En0 
    input [9:0] Pix_553, // sfix10_En0 
    input [9:0] Pix_554, // sfix10_En0 
    input [9:0] Pix_555, // sfix10_En0 
    input [9:0] Pix_556, // sfix10_En0 
    input [9:0] Pix_557, // sfix10_En0 
    input [9:0] Pix_558, // sfix10_En0 
    input [9:0] Pix_559, // sfix10_En0 
    input [9:0] Pix_560, // sfix10_En0 
    input [9:0] Pix_561, // sfix10_En0 
    input [9:0] Pix_562, // sfix10_En0 
    input [9:0] Pix_563, // sfix10_En0 
    input [9:0] Pix_564, // sfix10_En0 
    input [9:0] Pix_565, // sfix10_En0 
    input [9:0] Pix_566, // sfix10_En0 
    input [9:0] Pix_567, // sfix10_En0 
    input [9:0] Pix_568, // sfix10_En0 
    input [9:0] Pix_569, // sfix10_En0 
    input [9:0] Pix_570, // sfix10_En0 
    input [9:0] Pix_571, // sfix10_En0 
    input [9:0] Pix_572, // sfix10_En0 
    input [9:0] Pix_573, // sfix10_En0 
    input [9:0] Pix_574, // sfix10_En0 
    input [9:0] Pix_575, // sfix10_En0 
    input [9:0] Pix_576, // sfix10_En0 
    input [9:0] Pix_577, // sfix10_En0 
    input [9:0] Pix_578, // sfix10_En0 
    input [9:0] Pix_579, // sfix10_En0 
    input [9:0] Pix_580, // sfix10_En0 
    input [9:0] Pix_581, // sfix10_En0 
    input [9:0] Pix_582, // sfix10_En0 
    input [9:0] Pix_583, // sfix10_En0 
    input [9:0] Pix_584, // sfix10_En0 
    input [9:0] Pix_585, // sfix10_En0 
    input [9:0] Pix_586, // sfix10_En0 
    input [9:0] Pix_587, // sfix10_En0 
    input [9:0] Pix_588, // sfix10_En0 
    input [9:0] Pix_589, // sfix10_En0 
    input [9:0] Pix_590, // sfix10_En0 
    input [9:0] Pix_591, // sfix10_En0 
    input [9:0] Pix_592, // sfix10_En0 
    input [9:0] Pix_593, // sfix10_En0 
    input [9:0] Pix_594, // sfix10_En0 
    input [9:0] Pix_595, // sfix10_En0 
    input [9:0] Pix_596, // sfix10_En0 
    input [9:0] Pix_597, // sfix10_En0 
    input [9:0] Pix_598, // sfix10_En0 
    input [9:0] Pix_599, // sfix10_En0 
    input [9:0] Pix_600, // sfix10_En0 
    input [9:0] Pix_601, // sfix10_En0 
    input [9:0] Pix_602, // sfix10_En0 
    input [9:0] Pix_603, // sfix10_En0 
    input [9:0] Pix_604, // sfix10_En0 
    input [9:0] Pix_605, // sfix10_En0 
    input [9:0] Pix_606, // sfix10_En0 
    input [9:0] Pix_607, // sfix10_En0 
    input [9:0] Pix_608, // sfix10_En0 
    input [9:0] Pix_609, // sfix10_En0 
    input [9:0] Pix_610, // sfix10_En0 
    input [9:0] Pix_611, // sfix10_En0 
    input [9:0] Pix_612, // sfix10_En0 
    input [9:0] Pix_613, // sfix10_En0 
    input [9:0] Pix_614, // sfix10_En0 
    input [9:0] Pix_615, // sfix10_En0 
    input [9:0] Pix_616, // sfix10_En0 
    input [9:0] Pix_617, // sfix10_En0 
    input [9:0] Pix_618, // sfix10_En0 
    input [9:0] Pix_619, // sfix10_En0 
    input [9:0] Pix_620, // sfix10_En0 
    input [9:0] Pix_621, // sfix10_En0 
    input [9:0] Pix_622, // sfix10_En0 
    input [9:0] Pix_623, // sfix10_En0 
    input [9:0] Pix_624, // sfix10_En0 
    input [9:0] Pix_625, // sfix10_En0 
    input [9:0] Pix_626, // sfix10_En0 
    input [9:0] Pix_627, // sfix10_En0 
    input [9:0] Pix_628, // sfix10_En0 
    input [9:0] Pix_629, // sfix10_En0 
    input [9:0] Pix_630, // sfix10_En0 
    input [9:0] Pix_631, // sfix10_En0 
    input [9:0] Pix_632, // sfix10_En0 
    input [9:0] Pix_633, // sfix10_En0 
    input [9:0] Pix_634, // sfix10_En0 
    input [9:0] Pix_635, // sfix10_En0 
    input [9:0] Pix_636, // sfix10_En0 
    input [9:0] Pix_637, // sfix10_En0 
    input [9:0] Pix_638, // sfix10_En0 
    input [9:0] Pix_639, // sfix10_En0 
    input [9:0] Pix_640, // sfix10_En0 
    input [9:0] Pix_641, // sfix10_En0 
    input [9:0] Pix_642, // sfix10_En0 
    input [9:0] Pix_643, // sfix10_En0 
    input [9:0] Pix_644, // sfix10_En0 
    input [9:0] Pix_645, // sfix10_En0 
    input [9:0] Pix_646, // sfix10_En0 
    input [9:0] Pix_647, // sfix10_En0 
    input [9:0] Pix_648, // sfix10_En0 
    input [9:0] Pix_649, // sfix10_En0 
    input [9:0] Pix_650, // sfix10_En0 
    input [9:0] Pix_651, // sfix10_En0 
    input [9:0] Pix_652, // sfix10_En0 
    input [9:0] Pix_653, // sfix10_En0 
    input [9:0] Pix_654, // sfix10_En0 
    input [9:0] Pix_655, // sfix10_En0 
    input [9:0] Pix_656, // sfix10_En0 
    input [9:0] Pix_657, // sfix10_En0 
    input [9:0] Pix_658, // sfix10_En0 
    input [9:0] Pix_659, // sfix10_En0 
    input [9:0] Pix_660, // sfix10_En0 
    input [9:0] Pix_661, // sfix10_En0 
    input [9:0] Pix_662, // sfix10_En0 
    input [9:0] Pix_663, // sfix10_En0 
    input [9:0] Pix_664, // sfix10_En0 
    input [9:0] Pix_665, // sfix10_En0 
    input [9:0] Pix_666, // sfix10_En0 
    input [9:0] Pix_667, // sfix10_En0 
    input [9:0] Pix_668, // sfix10_En0 
    input [9:0] Pix_669, // sfix10_En0 
    input [9:0] Pix_670, // sfix10_En0 
    input [9:0] Pix_671, // sfix10_En0 
    input [9:0] Pix_672, // sfix10_En0 
    input [9:0] Pix_673, // sfix10_En0 
    input [9:0] Pix_674, // sfix10_En0 
    input [9:0] Pix_675, // sfix10_En0 
    input [9:0] Pix_676, // sfix10_En0 
    input [9:0] Pix_677, // sfix10_En0 
    input [9:0] Pix_678, // sfix10_En0 
    input [9:0] Pix_679, // sfix10_En0 
    input [9:0] Pix_680, // sfix10_En0 
    input [9:0] Pix_681, // sfix10_En0 
    input [9:0] Pix_682, // sfix10_En0 
    input [9:0] Pix_683, // sfix10_En0 
    input [9:0] Pix_684, // sfix10_En0 
    input [9:0] Pix_685, // sfix10_En0 
    input [9:0] Pix_686, // sfix10_En0 
    input [9:0] Pix_687, // sfix10_En0 
    input [9:0] Pix_688, // sfix10_En0 
    input [9:0] Pix_689, // sfix10_En0 
    input [9:0] Pix_690, // sfix10_En0 
    input [9:0] Pix_691, // sfix10_En0 
    input [9:0] Pix_692, // sfix10_En0 
    input [9:0] Pix_693, // sfix10_En0 
    input [9:0] Pix_694, // sfix10_En0 
    input [9:0] Pix_695, // sfix10_En0 
    input [9:0] Pix_696, // sfix10_En0 
    input [9:0] Pix_697, // sfix10_En0 
    input [9:0] Pix_698, // sfix10_En0 
    input [9:0] Pix_699, // sfix10_En0 
    input [9:0] Pix_700, // sfix10_En0 
    input [9:0] Pix_701, // sfix10_En0 
    input [9:0] Pix_702, // sfix10_En0 
    input [9:0] Pix_703, // sfix10_En0 
    input [9:0] Pix_704, // sfix10_En0 
    input [9:0] Pix_705, // sfix10_En0 
    input [9:0] Pix_706, // sfix10_En0 
    input [9:0] Pix_707, // sfix10_En0 
    input [9:0] Pix_708, // sfix10_En0 
    input [9:0] Pix_709, // sfix10_En0 
    input [9:0] Pix_710, // sfix10_En0 
    input [9:0] Pix_711, // sfix10_En0 
    input [9:0] Pix_712, // sfix10_En0 
    input [9:0] Pix_713, // sfix10_En0 
    input [9:0] Pix_714, // sfix10_En0 
    input [9:0] Pix_715, // sfix10_En0 
    input [9:0] Pix_716, // sfix10_En0 
    input [9:0] Pix_717, // sfix10_En0 
    input [9:0] Pix_718, // sfix10_En0 
    input [9:0] Pix_719, // sfix10_En0 
    input [9:0] Pix_720, // sfix10_En0 
    input [9:0] Pix_721, // sfix10_En0 
    input [9:0] Pix_722, // sfix10_En0 
    input [9:0] Pix_723, // sfix10_En0 
    input [9:0] Pix_724, // sfix10_En0 
    input [9:0] Pix_725, // sfix10_En0 
    input [9:0] Pix_726, // sfix10_En0 
    input [9:0] Pix_727, // sfix10_En0 
    input [9:0] Pix_728, // sfix10_En0 
    input [9:0] Pix_729, // sfix10_En0 
    input [9:0] Pix_730, // sfix10_En0 
    input [9:0] Pix_731, // sfix10_En0 
    input [9:0] Pix_732, // sfix10_En0 
    input [9:0] Pix_733, // sfix10_En0 
    input [9:0] Pix_734, // sfix10_En0 
    input [9:0] Pix_735, // sfix10_En0 
    input [9:0] Pix_736, // sfix10_En0 
    input [9:0] Pix_737, // sfix10_En0 
    input [9:0] Pix_738, // sfix10_En0 
    input [9:0] Pix_739, // sfix10_En0 
    input [9:0] Pix_740, // sfix10_En0 
    input [9:0] Pix_741, // sfix10_En0 
    input [9:0] Pix_742, // sfix10_En0 
    input [9:0] Pix_743, // sfix10_En0 
    input [9:0] Pix_744, // sfix10_En0 
    input [9:0] Pix_745, // sfix10_En0 
    input [9:0] Pix_746, // sfix10_En0 
    input [9:0] Pix_747, // sfix10_En0 
    input [9:0] Pix_748, // sfix10_En0 
    input [9:0] Pix_749, // sfix10_En0 
    input [9:0] Pix_750, // sfix10_En0 
    input [9:0] Pix_751, // sfix10_En0 
    input [9:0] Pix_752, // sfix10_En0 
    input [9:0] Pix_753, // sfix10_En0 
    input [9:0] Pix_754, // sfix10_En0 
    input [9:0] Pix_755, // sfix10_En0 
    input [9:0] Pix_756, // sfix10_En0 
    input [9:0] Pix_757, // sfix10_En0 
    input [9:0] Pix_758, // sfix10_En0 
    input [9:0] Pix_759, // sfix10_En0 
    input [9:0] Pix_760, // sfix10_En0 
    input [9:0] Pix_761, // sfix10_En0 
    input [9:0] Pix_762, // sfix10_En0 
    input [9:0] Pix_763, // sfix10_En0 
    input [9:0] Pix_764, // sfix10_En0 
    input [9:0] Pix_765, // sfix10_En0 
    input [9:0] Pix_766, // sfix10_En0 
    input [9:0] Pix_767, // sfix10_En0 
    input [9:0] Pix_768, // sfix10_En0 
    input [9:0] Pix_769, // sfix10_En0 
    input [9:0] Pix_770, // sfix10_En0 
    input [9:0] Pix_771, // sfix10_En0 
    input [9:0] Pix_772, // sfix10_En0 
    input [9:0] Pix_773, // sfix10_En0 
    input [9:0] Pix_774, // sfix10_En0 
    input [9:0] Pix_775, // sfix10_En0 
    input [9:0] Pix_776, // sfix10_En0 
    input [9:0] Pix_777, // sfix10_En0 
    input [9:0] Pix_778, // sfix10_En0 
    input [9:0] Pix_779, // sfix10_En0 
    input [9:0] Pix_780, // sfix10_En0 
    input [9:0] Pix_781, // sfix10_En0 
    input [9:0] Pix_782, // sfix10_En0 
    input [9:0] Pix_783, // sfix10_En0 
    input [9:0] Pix_784, // sfix10_En0 
 output [3:0] Image_Number, // sfix26_En18 
 output reg Output_Valid 
 );

//////// State Machine Formation////////
 reg[6:0] state, nxt_state;
 reg Load;
 always@(posedge clk, negedge GlobalReset) begin
     if(!GlobalReset) begin
        state <= 0;
     end
     else
        state <= nxt_state;
    end

//////// Regiser/Buffer Instanitaion////
// Buffers for max selecting
    reg[3:0] W11_n,W12_n,W13_n,W14_n,W15_n;
    reg signed[25:0] V11_n,V12_n,V13_n,V14_n,V15_n;
    reg[3:0] W21_n,W22_n;
    reg signed[25:0] V21_n,V22_n;
    reg[3:0] W31_n,W32_n;
    reg signed[25:0] V31_n,V32_n;

    reg[3:0] W11,W12,W13,W14,W15;
    reg signed[25:0] V11,V12,V13,V14,V15;
    reg[3:0] W21,W22;
    reg signed[25:0] V21,V22;
    reg[3:0] W31,W32;
    reg signed[25:0] V31,V32;
// Buffer for addition result
reg signed [25:0] Res0_n,Res1_n,Res2_n,Res3_n,Res4_n,Res5_n,Res6_n,Res7_n,Res8_n,Res9_n;
reg signed [25:0] Res0,Res1,Res2,Res3,Res4,Res5,Res6,Res7,Res8,Res9;
reg signed [25:0] Res_0_0,
    Res_0_1,
    Res_0_2,
    Res_0_3,
    Res_0_4,
    Res_0_5,
    Res_0_6,
    Res_0_7,
    Res_1_0,
    Res_1_1,
    Res_1_2,
    Res_1_3,
    Res_1_4,
    Res_1_5,
    Res_1_6,
    Res_1_7,
    Res_2_0,
    Res_2_1,
    Res_2_2,
    Res_2_3,
    Res_2_4,
    Res_2_5,
    Res_2_6,
    Res_2_7,
    Res_3_0,
    Res_3_1,
    Res_3_2,
    Res_3_3,
    Res_3_4,
    Res_3_5,
    Res_3_6,
    Res_3_7,
    Res_4_0,
    Res_4_1,
    Res_4_2,
    Res_4_3,
    Res_4_4,
    Res_4_5,
    Res_4_6,
    Res_4_7,
    Res_5_0,
    Res_5_1,
    Res_5_2,
    Res_5_3,
    Res_5_4,
    Res_5_5,
    Res_5_6,
    Res_5_7,
    Res_6_0,
    Res_6_1,
    Res_6_2,
    Res_6_3,
    Res_6_4,
    Res_6_5,
    Res_6_6,
    Res_6_7,
    Res_7_0,
    Res_7_1,
    Res_7_2,
    Res_7_3,
    Res_7_4,
    Res_7_5,
    Res_7_6,
    Res_7_7,
    Res_8_0,
    Res_8_1,
    Res_8_2,
    Res_8_3,
    Res_8_4,
    Res_8_5,
    Res_8_6,
    Res_8_7,
    Res_9_0,
    Res_9_1,
    Res_9_2,
    Res_9_3,
    Res_9_4,
    Res_9_5,
    Res_9_6,
    Res_9_7;

reg signed [25:0] Res_0_0_n,
    Res_0_1_n,
    Res_0_2_n,
    Res_0_3_n,
    Res_0_4_n,
    Res_0_5_n,
    Res_0_6_n,
    Res_0_7_n,
    Res_1_0_n,
    Res_1_1_n,
    Res_1_2_n,
    Res_1_3_n,
    Res_1_4_n,
    Res_1_5_n,
    Res_1_6_n,
    Res_1_7_n,
    Res_2_0_n,
    Res_2_1_n,
    Res_2_2_n,
    Res_2_3_n,
    Res_2_4_n,
    Res_2_5_n,
    Res_2_6_n,
    Res_2_7_n,
    Res_3_0_n,
    Res_3_1_n,
    Res_3_2_n,
    Res_3_3_n,
    Res_3_4_n,
    Res_3_5_n,
    Res_3_6_n,
    Res_3_7_n,
    Res_4_0_n,
    Res_4_1_n,
    Res_4_2_n,
    Res_4_3_n,
    Res_4_4_n,
    Res_4_5_n,
    Res_4_6_n,
    Res_4_7_n,
    Res_5_0_n,
    Res_5_1_n,
    Res_5_2_n,
    Res_5_3_n,
    Res_5_4_n,
    Res_5_5_n,
    Res_5_6_n,
    Res_5_7_n,
    Res_6_0_n,
    Res_6_1_n,
    Res_6_2_n,
    Res_6_3_n,
    Res_6_4_n,
    Res_6_5_n,
    Res_6_6_n,
    Res_6_7_n,
    Res_7_0_n,
    Res_7_1_n,
    Res_7_2_n,
    Res_7_3_n,
    Res_7_4_n,
    Res_7_5_n,
    Res_7_6_n,
    Res_7_7_n,
    Res_8_0_n,
    Res_8_1_n,
    Res_8_2_n,
    Res_8_3_n,
    Res_8_4_n,
    Res_8_5_n,
    Res_8_6_n,
    Res_8_7_n,
    Res_9_0_n,
    Res_9_1_n,
    Res_9_2_n,
    Res_9_3_n,
    Res_9_4_n,
    Res_9_5_n,
    Res_9_6_n,
    Res_9_7_n;
// Buffer for feature map input
reg[9:0] FeatureBuf_0;
    reg[9:0] FeatureBuf_1;
    reg[9:0] FeatureBuf_2;
    reg[9:0] FeatureBuf_3;
    reg[9:0] FeatureBuf_4;
    reg[9:0] FeatureBuf_5;
    reg[9:0] FeatureBuf_6;
    reg[9:0] FeatureBuf_7;
    reg[9:0] FeatureBuf_8;
    reg[9:0] FeatureBuf_9;
    reg[9:0] FeatureBuf_10;
    reg[9:0] FeatureBuf_11;
    reg[9:0] FeatureBuf_12;
    reg[9:0] FeatureBuf_13;
    reg[9:0] FeatureBuf_14;
    reg[9:0] FeatureBuf_15;
    reg[9:0] FeatureBuf_16;
    reg[9:0] FeatureBuf_17;
    reg[9:0] FeatureBuf_18;
    reg[9:0] FeatureBuf_19;
    reg[9:0] FeatureBuf_20;
    reg[9:0] FeatureBuf_21;
    reg[9:0] FeatureBuf_22;
    reg[9:0] FeatureBuf_23;
    reg[9:0] FeatureBuf_24;
    reg[9:0] FeatureBuf_25;
    reg[9:0] FeatureBuf_26;
    reg[9:0] FeatureBuf_27;
    reg[9:0] FeatureBuf_28;
    reg[9:0] FeatureBuf_29;
    reg[9:0] FeatureBuf_30;
    reg[9:0] FeatureBuf_31;
    reg[9:0] FeatureBuf_32;
    reg[9:0] FeatureBuf_33;
    reg[9:0] FeatureBuf_34;
    reg[9:0] FeatureBuf_35;
    reg[9:0] FeatureBuf_36;
    reg[9:0] FeatureBuf_37;
    reg[9:0] FeatureBuf_38;
    reg[9:0] FeatureBuf_39;
    reg[9:0] FeatureBuf_40;
    reg[9:0] FeatureBuf_41;
    reg[9:0] FeatureBuf_42;
    reg[9:0] FeatureBuf_43;
    reg[9:0] FeatureBuf_44;
    reg[9:0] FeatureBuf_45;
    reg[9:0] FeatureBuf_46;
    reg[9:0] FeatureBuf_47;
    reg[9:0] FeatureBuf_48;
    reg[9:0] FeatureBuf_49;
    reg[9:0] FeatureBuf_50;
    reg[9:0] FeatureBuf_51;
    reg[9:0] FeatureBuf_52;
    reg[9:0] FeatureBuf_53;
    reg[9:0] FeatureBuf_54;
    reg[9:0] FeatureBuf_55;
    reg[9:0] FeatureBuf_56;
    reg[9:0] FeatureBuf_57;
    reg[9:0] FeatureBuf_58;
    reg[9:0] FeatureBuf_59;
    reg[9:0] FeatureBuf_60;
    reg[9:0] FeatureBuf_61;
    reg[9:0] FeatureBuf_62;
    reg[9:0] FeatureBuf_63;
    reg[9:0] FeatureBuf_64;
    reg[9:0] FeatureBuf_65;
    reg[9:0] FeatureBuf_66;
    reg[9:0] FeatureBuf_67;
    reg[9:0] FeatureBuf_68;
    reg[9:0] FeatureBuf_69;
    reg[9:0] FeatureBuf_70;
    reg[9:0] FeatureBuf_71;
    reg[9:0] FeatureBuf_72;
    reg[9:0] FeatureBuf_73;
    reg[9:0] FeatureBuf_74;
    reg[9:0] FeatureBuf_75;
    reg[9:0] FeatureBuf_76;
    reg[9:0] FeatureBuf_77;
    reg[9:0] FeatureBuf_78;
    reg[9:0] FeatureBuf_79;
    reg[9:0] FeatureBuf_80;
    reg[9:0] FeatureBuf_81;
    reg[9:0] FeatureBuf_82;
    reg[9:0] FeatureBuf_83;
    reg[9:0] FeatureBuf_84;
    reg[9:0] FeatureBuf_85;
    reg[9:0] FeatureBuf_86;
    reg[9:0] FeatureBuf_87;
    reg[9:0] FeatureBuf_88;
    reg[9:0] FeatureBuf_89;
    reg[9:0] FeatureBuf_90;
    reg[9:0] FeatureBuf_91;
    reg[9:0] FeatureBuf_92;
    reg[9:0] FeatureBuf_93;
    reg[9:0] FeatureBuf_94;
    reg[9:0] FeatureBuf_95;
    reg[9:0] FeatureBuf_96;
    reg[9:0] FeatureBuf_97;
    reg[9:0] FeatureBuf_98;
    reg[9:0] FeatureBuf_99;
    reg[9:0] FeatureBuf_100;
    reg[9:0] FeatureBuf_101;
    reg[9:0] FeatureBuf_102;
    reg[9:0] FeatureBuf_103;
    reg[9:0] FeatureBuf_104;
    reg[9:0] FeatureBuf_105;
    reg[9:0] FeatureBuf_106;
    reg[9:0] FeatureBuf_107;
    reg[9:0] FeatureBuf_108;
    reg[9:0] FeatureBuf_109;
    reg[9:0] FeatureBuf_110;
    reg[9:0] FeatureBuf_111;
    reg[9:0] FeatureBuf_112;
    reg[9:0] FeatureBuf_113;
    reg[9:0] FeatureBuf_114;
    reg[9:0] FeatureBuf_115;
    reg[9:0] FeatureBuf_116;
    reg[9:0] FeatureBuf_117;
    reg[9:0] FeatureBuf_118;
    reg[9:0] FeatureBuf_119;
    reg[9:0] FeatureBuf_120;
    reg[9:0] FeatureBuf_121;
    reg[9:0] FeatureBuf_122;
    reg[9:0] FeatureBuf_123;
    reg[9:0] FeatureBuf_124;
    reg[9:0] FeatureBuf_125;
    reg[9:0] FeatureBuf_126;
    reg[9:0] FeatureBuf_127;
    reg[9:0] FeatureBuf_128;
    reg[9:0] FeatureBuf_129;
    reg[9:0] FeatureBuf_130;
    reg[9:0] FeatureBuf_131;
    reg[9:0] FeatureBuf_132;
    reg[9:0] FeatureBuf_133;
    reg[9:0] FeatureBuf_134;
    reg[9:0] FeatureBuf_135;
    reg[9:0] FeatureBuf_136;
    reg[9:0] FeatureBuf_137;
    reg[9:0] FeatureBuf_138;
    reg[9:0] FeatureBuf_139;
    reg[9:0] FeatureBuf_140;
    reg[9:0] FeatureBuf_141;
    reg[9:0] FeatureBuf_142;
    reg[9:0] FeatureBuf_143;
    reg[9:0] FeatureBuf_144;
    reg[9:0] FeatureBuf_145;
    reg[9:0] FeatureBuf_146;
    reg[9:0] FeatureBuf_147;
    reg[9:0] FeatureBuf_148;
    reg[9:0] FeatureBuf_149;
    reg[9:0] FeatureBuf_150;
    reg[9:0] FeatureBuf_151;
    reg[9:0] FeatureBuf_152;
    reg[9:0] FeatureBuf_153;
    reg[9:0] FeatureBuf_154;
    reg[9:0] FeatureBuf_155;
    reg[9:0] FeatureBuf_156;
    reg[9:0] FeatureBuf_157;
    reg[9:0] FeatureBuf_158;
    reg[9:0] FeatureBuf_159;
    reg[9:0] FeatureBuf_160;
    reg[9:0] FeatureBuf_161;
    reg[9:0] FeatureBuf_162;
    reg[9:0] FeatureBuf_163;
    reg[9:0] FeatureBuf_164;
    reg[9:0] FeatureBuf_165;
    reg[9:0] FeatureBuf_166;
    reg[9:0] FeatureBuf_167;
    reg[9:0] FeatureBuf_168;
    reg[9:0] FeatureBuf_169;
    reg[9:0] FeatureBuf_170;
    reg[9:0] FeatureBuf_171;
    reg[9:0] FeatureBuf_172;
    reg[9:0] FeatureBuf_173;
    reg[9:0] FeatureBuf_174;
    reg[9:0] FeatureBuf_175;
    reg[9:0] FeatureBuf_176;
    reg[9:0] FeatureBuf_177;
    reg[9:0] FeatureBuf_178;
    reg[9:0] FeatureBuf_179;
    reg[9:0] FeatureBuf_180;
    reg[9:0] FeatureBuf_181;
    reg[9:0] FeatureBuf_182;
    reg[9:0] FeatureBuf_183;
    reg[9:0] FeatureBuf_184;
    reg[9:0] FeatureBuf_185;
    reg[9:0] FeatureBuf_186;
    reg[9:0] FeatureBuf_187;
    reg[9:0] FeatureBuf_188;
    reg[9:0] FeatureBuf_189;
    reg[9:0] FeatureBuf_190;
    reg[9:0] FeatureBuf_191;
    reg[9:0] FeatureBuf_192;
    reg[9:0] FeatureBuf_193;
    reg[9:0] FeatureBuf_194;
    reg[9:0] FeatureBuf_195;
    reg[9:0] FeatureBuf_196;
    reg[9:0] FeatureBuf_197;
    reg[9:0] FeatureBuf_198;
    reg[9:0] FeatureBuf_199;
    reg[9:0] FeatureBuf_200;
    reg[9:0] FeatureBuf_201;
    reg[9:0] FeatureBuf_202;
    reg[9:0] FeatureBuf_203;
    reg[9:0] FeatureBuf_204;
    reg[9:0] FeatureBuf_205;
    reg[9:0] FeatureBuf_206;
    reg[9:0] FeatureBuf_207;
    reg[9:0] FeatureBuf_208;
    reg[9:0] FeatureBuf_209;
    reg[9:0] FeatureBuf_210;
    reg[9:0] FeatureBuf_211;
    reg[9:0] FeatureBuf_212;
    reg[9:0] FeatureBuf_213;
    reg[9:0] FeatureBuf_214;
    reg[9:0] FeatureBuf_215;
    reg[9:0] FeatureBuf_216;
    reg[9:0] FeatureBuf_217;
    reg[9:0] FeatureBuf_218;
    reg[9:0] FeatureBuf_219;
    reg[9:0] FeatureBuf_220;
    reg[9:0] FeatureBuf_221;
    reg[9:0] FeatureBuf_222;
    reg[9:0] FeatureBuf_223;
    reg[9:0] FeatureBuf_224;
    reg[9:0] FeatureBuf_225;
    reg[9:0] FeatureBuf_226;
    reg[9:0] FeatureBuf_227;
    reg[9:0] FeatureBuf_228;
    reg[9:0] FeatureBuf_229;
    reg[9:0] FeatureBuf_230;
    reg[9:0] FeatureBuf_231;
    reg[9:0] FeatureBuf_232;
    reg[9:0] FeatureBuf_233;
    reg[9:0] FeatureBuf_234;
    reg[9:0] FeatureBuf_235;
    reg[9:0] FeatureBuf_236;
    reg[9:0] FeatureBuf_237;
    reg[9:0] FeatureBuf_238;
    reg[9:0] FeatureBuf_239;
    reg[9:0] FeatureBuf_240;
    reg[9:0] FeatureBuf_241;
    reg[9:0] FeatureBuf_242;
    reg[9:0] FeatureBuf_243;
    reg[9:0] FeatureBuf_244;
    reg[9:0] FeatureBuf_245;
    reg[9:0] FeatureBuf_246;
    reg[9:0] FeatureBuf_247;
    reg[9:0] FeatureBuf_248;
    reg[9:0] FeatureBuf_249;
    reg[9:0] FeatureBuf_250;
    reg[9:0] FeatureBuf_251;
    reg[9:0] FeatureBuf_252;
    reg[9:0] FeatureBuf_253;
    reg[9:0] FeatureBuf_254;
    reg[9:0] FeatureBuf_255;
    reg[9:0] FeatureBuf_256;
    reg[9:0] FeatureBuf_257;
    reg[9:0] FeatureBuf_258;
    reg[9:0] FeatureBuf_259;
    reg[9:0] FeatureBuf_260;
    reg[9:0] FeatureBuf_261;
    reg[9:0] FeatureBuf_262;
    reg[9:0] FeatureBuf_263;
    reg[9:0] FeatureBuf_264;
    reg[9:0] FeatureBuf_265;
    reg[9:0] FeatureBuf_266;
    reg[9:0] FeatureBuf_267;
    reg[9:0] FeatureBuf_268;
    reg[9:0] FeatureBuf_269;
    reg[9:0] FeatureBuf_270;
    reg[9:0] FeatureBuf_271;
    reg[9:0] FeatureBuf_272;
    reg[9:0] FeatureBuf_273;
    reg[9:0] FeatureBuf_274;
    reg[9:0] FeatureBuf_275;
    reg[9:0] FeatureBuf_276;
    reg[9:0] FeatureBuf_277;
    reg[9:0] FeatureBuf_278;
    reg[9:0] FeatureBuf_279;
    reg[9:0] FeatureBuf_280;
    reg[9:0] FeatureBuf_281;
    reg[9:0] FeatureBuf_282;
    reg[9:0] FeatureBuf_283;
    reg[9:0] FeatureBuf_284;
    reg[9:0] FeatureBuf_285;
    reg[9:0] FeatureBuf_286;
    reg[9:0] FeatureBuf_287;
    reg[9:0] FeatureBuf_288;
    reg[9:0] FeatureBuf_289;
    reg[9:0] FeatureBuf_290;
    reg[9:0] FeatureBuf_291;
    reg[9:0] FeatureBuf_292;
    reg[9:0] FeatureBuf_293;
    reg[9:0] FeatureBuf_294;
    reg[9:0] FeatureBuf_295;
    reg[9:0] FeatureBuf_296;
    reg[9:0] FeatureBuf_297;
    reg[9:0] FeatureBuf_298;
    reg[9:0] FeatureBuf_299;
    reg[9:0] FeatureBuf_300;
    reg[9:0] FeatureBuf_301;
    reg[9:0] FeatureBuf_302;
    reg[9:0] FeatureBuf_303;
    reg[9:0] FeatureBuf_304;
    reg[9:0] FeatureBuf_305;
    reg[9:0] FeatureBuf_306;
    reg[9:0] FeatureBuf_307;
    reg[9:0] FeatureBuf_308;
    reg[9:0] FeatureBuf_309;
    reg[9:0] FeatureBuf_310;
    reg[9:0] FeatureBuf_311;
    reg[9:0] FeatureBuf_312;
    reg[9:0] FeatureBuf_313;
    reg[9:0] FeatureBuf_314;
    reg[9:0] FeatureBuf_315;
    reg[9:0] FeatureBuf_316;
    reg[9:0] FeatureBuf_317;
    reg[9:0] FeatureBuf_318;
    reg[9:0] FeatureBuf_319;
    reg[9:0] FeatureBuf_320;
    reg[9:0] FeatureBuf_321;
    reg[9:0] FeatureBuf_322;
    reg[9:0] FeatureBuf_323;
    reg[9:0] FeatureBuf_324;
    reg[9:0] FeatureBuf_325;
    reg[9:0] FeatureBuf_326;
    reg[9:0] FeatureBuf_327;
    reg[9:0] FeatureBuf_328;
    reg[9:0] FeatureBuf_329;
    reg[9:0] FeatureBuf_330;
    reg[9:0] FeatureBuf_331;
    reg[9:0] FeatureBuf_332;
    reg[9:0] FeatureBuf_333;
    reg[9:0] FeatureBuf_334;
    reg[9:0] FeatureBuf_335;
    reg[9:0] FeatureBuf_336;
    reg[9:0] FeatureBuf_337;
    reg[9:0] FeatureBuf_338;
    reg[9:0] FeatureBuf_339;
    reg[9:0] FeatureBuf_340;
    reg[9:0] FeatureBuf_341;
    reg[9:0] FeatureBuf_342;
    reg[9:0] FeatureBuf_343;
    reg[9:0] FeatureBuf_344;
    reg[9:0] FeatureBuf_345;
    reg[9:0] FeatureBuf_346;
    reg[9:0] FeatureBuf_347;
    reg[9:0] FeatureBuf_348;
    reg[9:0] FeatureBuf_349;
    reg[9:0] FeatureBuf_350;
    reg[9:0] FeatureBuf_351;
    reg[9:0] FeatureBuf_352;
    reg[9:0] FeatureBuf_353;
    reg[9:0] FeatureBuf_354;
    reg[9:0] FeatureBuf_355;
    reg[9:0] FeatureBuf_356;
    reg[9:0] FeatureBuf_357;
    reg[9:0] FeatureBuf_358;
    reg[9:0] FeatureBuf_359;
    reg[9:0] FeatureBuf_360;
    reg[9:0] FeatureBuf_361;
    reg[9:0] FeatureBuf_362;
    reg[9:0] FeatureBuf_363;
    reg[9:0] FeatureBuf_364;
    reg[9:0] FeatureBuf_365;
    reg[9:0] FeatureBuf_366;
    reg[9:0] FeatureBuf_367;
    reg[9:0] FeatureBuf_368;
    reg[9:0] FeatureBuf_369;
    reg[9:0] FeatureBuf_370;
    reg[9:0] FeatureBuf_371;
    reg[9:0] FeatureBuf_372;
    reg[9:0] FeatureBuf_373;
    reg[9:0] FeatureBuf_374;
    reg[9:0] FeatureBuf_375;
    reg[9:0] FeatureBuf_376;
    reg[9:0] FeatureBuf_377;
    reg[9:0] FeatureBuf_378;
    reg[9:0] FeatureBuf_379;
    reg[9:0] FeatureBuf_380;
    reg[9:0] FeatureBuf_381;
    reg[9:0] FeatureBuf_382;
    reg[9:0] FeatureBuf_383;
    reg[9:0] FeatureBuf_384;
    reg[9:0] FeatureBuf_385;
    reg[9:0] FeatureBuf_386;
    reg[9:0] FeatureBuf_387;
    reg[9:0] FeatureBuf_388;
    reg[9:0] FeatureBuf_389;
    reg[9:0] FeatureBuf_390;
    reg[9:0] FeatureBuf_391;
    reg[9:0] FeatureBuf_392;
    reg[9:0] FeatureBuf_393;
    reg[9:0] FeatureBuf_394;
    reg[9:0] FeatureBuf_395;
    reg[9:0] FeatureBuf_396;
    reg[9:0] FeatureBuf_397;
    reg[9:0] FeatureBuf_398;
    reg[9:0] FeatureBuf_399;
    reg[9:0] FeatureBuf_400;
    reg[9:0] FeatureBuf_401;
    reg[9:0] FeatureBuf_402;
    reg[9:0] FeatureBuf_403;
    reg[9:0] FeatureBuf_404;
    reg[9:0] FeatureBuf_405;
    reg[9:0] FeatureBuf_406;
    reg[9:0] FeatureBuf_407;
    reg[9:0] FeatureBuf_408;
    reg[9:0] FeatureBuf_409;
    reg[9:0] FeatureBuf_410;
    reg[9:0] FeatureBuf_411;
    reg[9:0] FeatureBuf_412;
    reg[9:0] FeatureBuf_413;
    reg[9:0] FeatureBuf_414;
    reg[9:0] FeatureBuf_415;
    reg[9:0] FeatureBuf_416;
    reg[9:0] FeatureBuf_417;
    reg[9:0] FeatureBuf_418;
    reg[9:0] FeatureBuf_419;
    reg[9:0] FeatureBuf_420;
    reg[9:0] FeatureBuf_421;
    reg[9:0] FeatureBuf_422;
    reg[9:0] FeatureBuf_423;
    reg[9:0] FeatureBuf_424;
    reg[9:0] FeatureBuf_425;
    reg[9:0] FeatureBuf_426;
    reg[9:0] FeatureBuf_427;
    reg[9:0] FeatureBuf_428;
    reg[9:0] FeatureBuf_429;
    reg[9:0] FeatureBuf_430;
    reg[9:0] FeatureBuf_431;
    reg[9:0] FeatureBuf_432;
    reg[9:0] FeatureBuf_433;
    reg[9:0] FeatureBuf_434;
    reg[9:0] FeatureBuf_435;
    reg[9:0] FeatureBuf_436;
    reg[9:0] FeatureBuf_437;
    reg[9:0] FeatureBuf_438;
    reg[9:0] FeatureBuf_439;
    reg[9:0] FeatureBuf_440;
    reg[9:0] FeatureBuf_441;
    reg[9:0] FeatureBuf_442;
    reg[9:0] FeatureBuf_443;
    reg[9:0] FeatureBuf_444;
    reg[9:0] FeatureBuf_445;
    reg[9:0] FeatureBuf_446;
    reg[9:0] FeatureBuf_447;
    reg[9:0] FeatureBuf_448;
    reg[9:0] FeatureBuf_449;
    reg[9:0] FeatureBuf_450;
    reg[9:0] FeatureBuf_451;
    reg[9:0] FeatureBuf_452;
    reg[9:0] FeatureBuf_453;
    reg[9:0] FeatureBuf_454;
    reg[9:0] FeatureBuf_455;
    reg[9:0] FeatureBuf_456;
    reg[9:0] FeatureBuf_457;
    reg[9:0] FeatureBuf_458;
    reg[9:0] FeatureBuf_459;
    reg[9:0] FeatureBuf_460;
    reg[9:0] FeatureBuf_461;
    reg[9:0] FeatureBuf_462;
    reg[9:0] FeatureBuf_463;
    reg[9:0] FeatureBuf_464;
    reg[9:0] FeatureBuf_465;
    reg[9:0] FeatureBuf_466;
    reg[9:0] FeatureBuf_467;
    reg[9:0] FeatureBuf_468;
    reg[9:0] FeatureBuf_469;
    reg[9:0] FeatureBuf_470;
    reg[9:0] FeatureBuf_471;
    reg[9:0] FeatureBuf_472;
    reg[9:0] FeatureBuf_473;
    reg[9:0] FeatureBuf_474;
    reg[9:0] FeatureBuf_475;
    reg[9:0] FeatureBuf_476;
    reg[9:0] FeatureBuf_477;
    reg[9:0] FeatureBuf_478;
    reg[9:0] FeatureBuf_479;
    reg[9:0] FeatureBuf_480;
    reg[9:0] FeatureBuf_481;
    reg[9:0] FeatureBuf_482;
    reg[9:0] FeatureBuf_483;
    reg[9:0] FeatureBuf_484;
    reg[9:0] FeatureBuf_485;
    reg[9:0] FeatureBuf_486;
    reg[9:0] FeatureBuf_487;
    reg[9:0] FeatureBuf_488;
    reg[9:0] FeatureBuf_489;
    reg[9:0] FeatureBuf_490;
    reg[9:0] FeatureBuf_491;
    reg[9:0] FeatureBuf_492;
    reg[9:0] FeatureBuf_493;
    reg[9:0] FeatureBuf_494;
    reg[9:0] FeatureBuf_495;
    reg[9:0] FeatureBuf_496;
    reg[9:0] FeatureBuf_497;
    reg[9:0] FeatureBuf_498;
    reg[9:0] FeatureBuf_499;
    reg[9:0] FeatureBuf_500;
    reg[9:0] FeatureBuf_501;
    reg[9:0] FeatureBuf_502;
    reg[9:0] FeatureBuf_503;
    reg[9:0] FeatureBuf_504;
    reg[9:0] FeatureBuf_505;
    reg[9:0] FeatureBuf_506;
    reg[9:0] FeatureBuf_507;
    reg[9:0] FeatureBuf_508;
    reg[9:0] FeatureBuf_509;
    reg[9:0] FeatureBuf_510;
    reg[9:0] FeatureBuf_511;
    reg[9:0] FeatureBuf_512;
    reg[9:0] FeatureBuf_513;
    reg[9:0] FeatureBuf_514;
    reg[9:0] FeatureBuf_515;
    reg[9:0] FeatureBuf_516;
    reg[9:0] FeatureBuf_517;
    reg[9:0] FeatureBuf_518;
    reg[9:0] FeatureBuf_519;
    reg[9:0] FeatureBuf_520;
    reg[9:0] FeatureBuf_521;
    reg[9:0] FeatureBuf_522;
    reg[9:0] FeatureBuf_523;
    reg[9:0] FeatureBuf_524;
    reg[9:0] FeatureBuf_525;
    reg[9:0] FeatureBuf_526;
    reg[9:0] FeatureBuf_527;
    reg[9:0] FeatureBuf_528;
    reg[9:0] FeatureBuf_529;
    reg[9:0] FeatureBuf_530;
    reg[9:0] FeatureBuf_531;
    reg[9:0] FeatureBuf_532;
    reg[9:0] FeatureBuf_533;
    reg[9:0] FeatureBuf_534;
    reg[9:0] FeatureBuf_535;
    reg[9:0] FeatureBuf_536;
    reg[9:0] FeatureBuf_537;
    reg[9:0] FeatureBuf_538;
    reg[9:0] FeatureBuf_539;
    reg[9:0] FeatureBuf_540;
    reg[9:0] FeatureBuf_541;
    reg[9:0] FeatureBuf_542;
    reg[9:0] FeatureBuf_543;
    reg[9:0] FeatureBuf_544;
    reg[9:0] FeatureBuf_545;
    reg[9:0] FeatureBuf_546;
    reg[9:0] FeatureBuf_547;
    reg[9:0] FeatureBuf_548;
    reg[9:0] FeatureBuf_549;
    reg[9:0] FeatureBuf_550;
    reg[9:0] FeatureBuf_551;
    reg[9:0] FeatureBuf_552;
    reg[9:0] FeatureBuf_553;
    reg[9:0] FeatureBuf_554;
    reg[9:0] FeatureBuf_555;
    reg[9:0] FeatureBuf_556;
    reg[9:0] FeatureBuf_557;
    reg[9:0] FeatureBuf_558;
    reg[9:0] FeatureBuf_559;
    reg[9:0] FeatureBuf_560;
    reg[9:0] FeatureBuf_561;
    reg[9:0] FeatureBuf_562;
    reg[9:0] FeatureBuf_563;
    reg[9:0] FeatureBuf_564;
    reg[9:0] FeatureBuf_565;
    reg[9:0] FeatureBuf_566;
    reg[9:0] FeatureBuf_567;
    reg[9:0] FeatureBuf_568;
    reg[9:0] FeatureBuf_569;
    reg[9:0] FeatureBuf_570;
    reg[9:0] FeatureBuf_571;
    reg[9:0] FeatureBuf_572;
    reg[9:0] FeatureBuf_573;
    reg[9:0] FeatureBuf_574;
    reg[9:0] FeatureBuf_575;
    reg[9:0] FeatureBuf_576;
    reg[9:0] FeatureBuf_577;
    reg[9:0] FeatureBuf_578;
    reg[9:0] FeatureBuf_579;
    reg[9:0] FeatureBuf_580;
    reg[9:0] FeatureBuf_581;
    reg[9:0] FeatureBuf_582;
    reg[9:0] FeatureBuf_583;
    reg[9:0] FeatureBuf_584;
    reg[9:0] FeatureBuf_585;
    reg[9:0] FeatureBuf_586;
    reg[9:0] FeatureBuf_587;
    reg[9:0] FeatureBuf_588;
    reg[9:0] FeatureBuf_589;
    reg[9:0] FeatureBuf_590;
    reg[9:0] FeatureBuf_591;
    reg[9:0] FeatureBuf_592;
    reg[9:0] FeatureBuf_593;
    reg[9:0] FeatureBuf_594;
    reg[9:0] FeatureBuf_595;
    reg[9:0] FeatureBuf_596;
    reg[9:0] FeatureBuf_597;
    reg[9:0] FeatureBuf_598;
    reg[9:0] FeatureBuf_599;
    reg[9:0] FeatureBuf_600;
    reg[9:0] FeatureBuf_601;
    reg[9:0] FeatureBuf_602;
    reg[9:0] FeatureBuf_603;
    reg[9:0] FeatureBuf_604;
    reg[9:0] FeatureBuf_605;
    reg[9:0] FeatureBuf_606;
    reg[9:0] FeatureBuf_607;
    reg[9:0] FeatureBuf_608;
    reg[9:0] FeatureBuf_609;
    reg[9:0] FeatureBuf_610;
    reg[9:0] FeatureBuf_611;
    reg[9:0] FeatureBuf_612;
    reg[9:0] FeatureBuf_613;
    reg[9:0] FeatureBuf_614;
    reg[9:0] FeatureBuf_615;
    reg[9:0] FeatureBuf_616;
    reg[9:0] FeatureBuf_617;
    reg[9:0] FeatureBuf_618;
    reg[9:0] FeatureBuf_619;
    reg[9:0] FeatureBuf_620;
    reg[9:0] FeatureBuf_621;
    reg[9:0] FeatureBuf_622;
    reg[9:0] FeatureBuf_623;
    reg[9:0] FeatureBuf_624;
    reg[9:0] FeatureBuf_625;
    reg[9:0] FeatureBuf_626;
    reg[9:0] FeatureBuf_627;
    reg[9:0] FeatureBuf_628;
    reg[9:0] FeatureBuf_629;
    reg[9:0] FeatureBuf_630;
    reg[9:0] FeatureBuf_631;
    reg[9:0] FeatureBuf_632;
    reg[9:0] FeatureBuf_633;
    reg[9:0] FeatureBuf_634;
    reg[9:0] FeatureBuf_635;
    reg[9:0] FeatureBuf_636;
    reg[9:0] FeatureBuf_637;
    reg[9:0] FeatureBuf_638;
    reg[9:0] FeatureBuf_639;
    reg[9:0] FeatureBuf_640;
    reg[9:0] FeatureBuf_641;
    reg[9:0] FeatureBuf_642;
    reg[9:0] FeatureBuf_643;
    reg[9:0] FeatureBuf_644;
    reg[9:0] FeatureBuf_645;
    reg[9:0] FeatureBuf_646;
    reg[9:0] FeatureBuf_647;
    reg[9:0] FeatureBuf_648;
    reg[9:0] FeatureBuf_649;
    reg[9:0] FeatureBuf_650;
    reg[9:0] FeatureBuf_651;
    reg[9:0] FeatureBuf_652;
    reg[9:0] FeatureBuf_653;
    reg[9:0] FeatureBuf_654;
    reg[9:0] FeatureBuf_655;
    reg[9:0] FeatureBuf_656;
    reg[9:0] FeatureBuf_657;
    reg[9:0] FeatureBuf_658;
    reg[9:0] FeatureBuf_659;
    reg[9:0] FeatureBuf_660;
    reg[9:0] FeatureBuf_661;
    reg[9:0] FeatureBuf_662;
    reg[9:0] FeatureBuf_663;
    reg[9:0] FeatureBuf_664;
    reg[9:0] FeatureBuf_665;
    reg[9:0] FeatureBuf_666;
    reg[9:0] FeatureBuf_667;
    reg[9:0] FeatureBuf_668;
    reg[9:0] FeatureBuf_669;
    reg[9:0] FeatureBuf_670;
    reg[9:0] FeatureBuf_671;
    reg[9:0] FeatureBuf_672;
    reg[9:0] FeatureBuf_673;
    reg[9:0] FeatureBuf_674;
    reg[9:0] FeatureBuf_675;
    reg[9:0] FeatureBuf_676;
    reg[9:0] FeatureBuf_677;
    reg[9:0] FeatureBuf_678;
    reg[9:0] FeatureBuf_679;
    reg[9:0] FeatureBuf_680;
    reg[9:0] FeatureBuf_681;
    reg[9:0] FeatureBuf_682;
    reg[9:0] FeatureBuf_683;
    reg[9:0] FeatureBuf_684;
    reg[9:0] FeatureBuf_685;
    reg[9:0] FeatureBuf_686;
    reg[9:0] FeatureBuf_687;
    reg[9:0] FeatureBuf_688;
    reg[9:0] FeatureBuf_689;
    reg[9:0] FeatureBuf_690;
    reg[9:0] FeatureBuf_691;
    reg[9:0] FeatureBuf_692;
    reg[9:0] FeatureBuf_693;
    reg[9:0] FeatureBuf_694;
    reg[9:0] FeatureBuf_695;
    reg[9:0] FeatureBuf_696;
    reg[9:0] FeatureBuf_697;
    reg[9:0] FeatureBuf_698;
    reg[9:0] FeatureBuf_699;
    reg[9:0] FeatureBuf_700;
    reg[9:0] FeatureBuf_701;
    reg[9:0] FeatureBuf_702;
    reg[9:0] FeatureBuf_703;
    reg[9:0] FeatureBuf_704;
    reg[9:0] FeatureBuf_705;
    reg[9:0] FeatureBuf_706;
    reg[9:0] FeatureBuf_707;
    reg[9:0] FeatureBuf_708;
    reg[9:0] FeatureBuf_709;
    reg[9:0] FeatureBuf_710;
    reg[9:0] FeatureBuf_711;
    reg[9:0] FeatureBuf_712;
    reg[9:0] FeatureBuf_713;
    reg[9:0] FeatureBuf_714;
    reg[9:0] FeatureBuf_715;
    reg[9:0] FeatureBuf_716;
    reg[9:0] FeatureBuf_717;
    reg[9:0] FeatureBuf_718;
    reg[9:0] FeatureBuf_719;
    reg[9:0] FeatureBuf_720;
    reg[9:0] FeatureBuf_721;
    reg[9:0] FeatureBuf_722;
    reg[9:0] FeatureBuf_723;
    reg[9:0] FeatureBuf_724;
    reg[9:0] FeatureBuf_725;
    reg[9:0] FeatureBuf_726;
    reg[9:0] FeatureBuf_727;
    reg[9:0] FeatureBuf_728;
    reg[9:0] FeatureBuf_729;
    reg[9:0] FeatureBuf_730;
    reg[9:0] FeatureBuf_731;
    reg[9:0] FeatureBuf_732;
    reg[9:0] FeatureBuf_733;
    reg[9:0] FeatureBuf_734;
    reg[9:0] FeatureBuf_735;
    reg[9:0] FeatureBuf_736;
    reg[9:0] FeatureBuf_737;
    reg[9:0] FeatureBuf_738;
    reg[9:0] FeatureBuf_739;
    reg[9:0] FeatureBuf_740;
    reg[9:0] FeatureBuf_741;
    reg[9:0] FeatureBuf_742;
    reg[9:0] FeatureBuf_743;
    reg[9:0] FeatureBuf_744;
    reg[9:0] FeatureBuf_745;
    reg[9:0] FeatureBuf_746;
    reg[9:0] FeatureBuf_747;
    reg[9:0] FeatureBuf_748;
    reg[9:0] FeatureBuf_749;
    reg[9:0] FeatureBuf_750;
    reg[9:0] FeatureBuf_751;
    reg[9:0] FeatureBuf_752;
    reg[9:0] FeatureBuf_753;
    reg[9:0] FeatureBuf_754;
    reg[9:0] FeatureBuf_755;
    reg[9:0] FeatureBuf_756;
    reg[9:0] FeatureBuf_757;
    reg[9:0] FeatureBuf_758;
    reg[9:0] FeatureBuf_759;
    reg[9:0] FeatureBuf_760;
    reg[9:0] FeatureBuf_761;
    reg[9:0] FeatureBuf_762;
    reg[9:0] FeatureBuf_763;
    reg[9:0] FeatureBuf_764;
    reg[9:0] FeatureBuf_765;
    reg[9:0] FeatureBuf_766;
    reg[9:0] FeatureBuf_767;
    reg[9:0] FeatureBuf_768;
    reg[9:0] FeatureBuf_769;
    reg[9:0] FeatureBuf_770;
    reg[9:0] FeatureBuf_771;
    reg[9:0] FeatureBuf_772;
    reg[9:0] FeatureBuf_773;
    reg[9:0] FeatureBuf_774;
    reg[9:0] FeatureBuf_775;
    reg[9:0] FeatureBuf_776;
    reg[9:0] FeatureBuf_777;
    reg[9:0] FeatureBuf_778;
    reg[9:0] FeatureBuf_779;
    reg[9:0] FeatureBuf_780;
    reg[9:0] FeatureBuf_781;
    reg[9:0] FeatureBuf_782;
    reg[9:0] FeatureBuf_783;

always@(posedge clk, negedge GlobalReset)begin
    if(!GlobalReset)begin
        W11 <= 0;
        W12 <= 0;
        W13 <= 0;
        W14 <= 0;
        W15 <= 0;
        V11 <= 0;
        V12 <= 0;
        V13 <= 0;
        V14 <= 0;
        V15 <= 0;
        W21 <= 0;
        W22 <= 0;
        V21 <= 0;
        V22 <= 0;
        W31 <= 0;
        W32 <= 0;
        V31 <= 0;
        V32 <= 0;
    end
    else  begin
        W11 <= W11_n;
        W12 <= W12_n;
        W13 <= W13_n;
        W14 <= W14_n;
        W15 <= W15_n;
        V11 <= V11_n;
        V12 <= V12_n;
        V13 <= V13_n;
        V14 <= V14_n;
        V15 <= V15_n;
        W21 <= W21_n;
        W22 <= W22_n;
        V21 <= V21_n;
        V22 <= V22_n;
        W31 <= W31_n;
        W32 <= W32_n;
        V31 <= V31_n;
        V32 <= V32_n;
    end
end

always@(posedge clk, negedge GlobalReset)begin
    if(!GlobalReset)begin
        FeatureBuf_0 <= 0;
        FeatureBuf_1 <= 0;
        FeatureBuf_2 <= 0;
        FeatureBuf_3 <= 0;
        FeatureBuf_4 <= 0;
        FeatureBuf_5 <= 0;
        FeatureBuf_6 <= 0;
        FeatureBuf_7 <= 0;
        FeatureBuf_8 <= 0;
        FeatureBuf_9 <= 0;
        FeatureBuf_10 <= 0;
        FeatureBuf_11 <= 0;
        FeatureBuf_12 <= 0;
        FeatureBuf_13 <= 0;
        FeatureBuf_14 <= 0;
        FeatureBuf_15 <= 0;
        FeatureBuf_16 <= 0;
        FeatureBuf_17 <= 0;
        FeatureBuf_18 <= 0;
        FeatureBuf_19 <= 0;
        FeatureBuf_20 <= 0;
        FeatureBuf_21 <= 0;
        FeatureBuf_22 <= 0;
        FeatureBuf_23 <= 0;
        FeatureBuf_24 <= 0;
        FeatureBuf_25 <= 0;
        FeatureBuf_26 <= 0;
        FeatureBuf_27 <= 0;
        FeatureBuf_28 <= 0;
        FeatureBuf_29 <= 0;
        FeatureBuf_30 <= 0;
        FeatureBuf_31 <= 0;
        FeatureBuf_32 <= 0;
        FeatureBuf_33 <= 0;
        FeatureBuf_34 <= 0;
        FeatureBuf_35 <= 0;
        FeatureBuf_36 <= 0;
        FeatureBuf_37 <= 0;
        FeatureBuf_38 <= 0;
        FeatureBuf_39 <= 0;
        FeatureBuf_40 <= 0;
        FeatureBuf_41 <= 0;
        FeatureBuf_42 <= 0;
        FeatureBuf_43 <= 0;
        FeatureBuf_44 <= 0;
        FeatureBuf_45 <= 0;
        FeatureBuf_46 <= 0;
        FeatureBuf_47 <= 0;
        FeatureBuf_48 <= 0;
        FeatureBuf_49 <= 0;
        FeatureBuf_50 <= 0;
        FeatureBuf_51 <= 0;
        FeatureBuf_52 <= 0;
        FeatureBuf_53 <= 0;
        FeatureBuf_54 <= 0;
        FeatureBuf_55 <= 0;
        FeatureBuf_56 <= 0;
        FeatureBuf_57 <= 0;
        FeatureBuf_58 <= 0;
        FeatureBuf_59 <= 0;
        FeatureBuf_60 <= 0;
        FeatureBuf_61 <= 0;
        FeatureBuf_62 <= 0;
        FeatureBuf_63 <= 0;
        FeatureBuf_64 <= 0;
        FeatureBuf_65 <= 0;
        FeatureBuf_66 <= 0;
        FeatureBuf_67 <= 0;
        FeatureBuf_68 <= 0;
        FeatureBuf_69 <= 0;
        FeatureBuf_70 <= 0;
        FeatureBuf_71 <= 0;
        FeatureBuf_72 <= 0;
        FeatureBuf_73 <= 0;
        FeatureBuf_74 <= 0;
        FeatureBuf_75 <= 0;
        FeatureBuf_76 <= 0;
        FeatureBuf_77 <= 0;
        FeatureBuf_78 <= 0;
        FeatureBuf_79 <= 0;
        FeatureBuf_80 <= 0;
        FeatureBuf_81 <= 0;
        FeatureBuf_82 <= 0;
        FeatureBuf_83 <= 0;
        FeatureBuf_84 <= 0;
        FeatureBuf_85 <= 0;
        FeatureBuf_86 <= 0;
        FeatureBuf_87 <= 0;
        FeatureBuf_88 <= 0;
        FeatureBuf_89 <= 0;
        FeatureBuf_90 <= 0;
        FeatureBuf_91 <= 0;
        FeatureBuf_92 <= 0;
        FeatureBuf_93 <= 0;
        FeatureBuf_94 <= 0;
        FeatureBuf_95 <= 0;
        FeatureBuf_96 <= 0;
        FeatureBuf_97 <= 0;
        FeatureBuf_98 <= 0;
        FeatureBuf_99 <= 0;
        FeatureBuf_100 <= 0;
        FeatureBuf_101 <= 0;
        FeatureBuf_102 <= 0;
        FeatureBuf_103 <= 0;
        FeatureBuf_104 <= 0;
        FeatureBuf_105 <= 0;
        FeatureBuf_106 <= 0;
        FeatureBuf_107 <= 0;
        FeatureBuf_108 <= 0;
        FeatureBuf_109 <= 0;
        FeatureBuf_110 <= 0;
        FeatureBuf_111 <= 0;
        FeatureBuf_112 <= 0;
        FeatureBuf_113 <= 0;
        FeatureBuf_114 <= 0;
        FeatureBuf_115 <= 0;
        FeatureBuf_116 <= 0;
        FeatureBuf_117 <= 0;
        FeatureBuf_118 <= 0;
        FeatureBuf_119 <= 0;
        FeatureBuf_120 <= 0;
        FeatureBuf_121 <= 0;
        FeatureBuf_122 <= 0;
        FeatureBuf_123 <= 0;
        FeatureBuf_124 <= 0;
        FeatureBuf_125 <= 0;
        FeatureBuf_126 <= 0;
        FeatureBuf_127 <= 0;
        FeatureBuf_128 <= 0;
        FeatureBuf_129 <= 0;
        FeatureBuf_130 <= 0;
        FeatureBuf_131 <= 0;
        FeatureBuf_132 <= 0;
        FeatureBuf_133 <= 0;
        FeatureBuf_134 <= 0;
        FeatureBuf_135 <= 0;
        FeatureBuf_136 <= 0;
        FeatureBuf_137 <= 0;
        FeatureBuf_138 <= 0;
        FeatureBuf_139 <= 0;
        FeatureBuf_140 <= 0;
        FeatureBuf_141 <= 0;
        FeatureBuf_142 <= 0;
        FeatureBuf_143 <= 0;
        FeatureBuf_144 <= 0;
        FeatureBuf_145 <= 0;
        FeatureBuf_146 <= 0;
        FeatureBuf_147 <= 0;
        FeatureBuf_148 <= 0;
        FeatureBuf_149 <= 0;
        FeatureBuf_150 <= 0;
        FeatureBuf_151 <= 0;
        FeatureBuf_152 <= 0;
        FeatureBuf_153 <= 0;
        FeatureBuf_154 <= 0;
        FeatureBuf_155 <= 0;
        FeatureBuf_156 <= 0;
        FeatureBuf_157 <= 0;
        FeatureBuf_158 <= 0;
        FeatureBuf_159 <= 0;
        FeatureBuf_160 <= 0;
        FeatureBuf_161 <= 0;
        FeatureBuf_162 <= 0;
        FeatureBuf_163 <= 0;
        FeatureBuf_164 <= 0;
        FeatureBuf_165 <= 0;
        FeatureBuf_166 <= 0;
        FeatureBuf_167 <= 0;
        FeatureBuf_168 <= 0;
        FeatureBuf_169 <= 0;
        FeatureBuf_170 <= 0;
        FeatureBuf_171 <= 0;
        FeatureBuf_172 <= 0;
        FeatureBuf_173 <= 0;
        FeatureBuf_174 <= 0;
        FeatureBuf_175 <= 0;
        FeatureBuf_176 <= 0;
        FeatureBuf_177 <= 0;
        FeatureBuf_178 <= 0;
        FeatureBuf_179 <= 0;
        FeatureBuf_180 <= 0;
        FeatureBuf_181 <= 0;
        FeatureBuf_182 <= 0;
        FeatureBuf_183 <= 0;
        FeatureBuf_184 <= 0;
        FeatureBuf_185 <= 0;
        FeatureBuf_186 <= 0;
        FeatureBuf_187 <= 0;
        FeatureBuf_188 <= 0;
        FeatureBuf_189 <= 0;
        FeatureBuf_190 <= 0;
        FeatureBuf_191 <= 0;
        FeatureBuf_192 <= 0;
        FeatureBuf_193 <= 0;
        FeatureBuf_194 <= 0;
        FeatureBuf_195 <= 0;
        FeatureBuf_196 <= 0;
        FeatureBuf_197 <= 0;
        FeatureBuf_198 <= 0;
        FeatureBuf_199 <= 0;
        FeatureBuf_200 <= 0;
        FeatureBuf_201 <= 0;
        FeatureBuf_202 <= 0;
        FeatureBuf_203 <= 0;
        FeatureBuf_204 <= 0;
        FeatureBuf_205 <= 0;
        FeatureBuf_206 <= 0;
        FeatureBuf_207 <= 0;
        FeatureBuf_208 <= 0;
        FeatureBuf_209 <= 0;
        FeatureBuf_210 <= 0;
        FeatureBuf_211 <= 0;
        FeatureBuf_212 <= 0;
        FeatureBuf_213 <= 0;
        FeatureBuf_214 <= 0;
        FeatureBuf_215 <= 0;
        FeatureBuf_216 <= 0;
        FeatureBuf_217 <= 0;
        FeatureBuf_218 <= 0;
        FeatureBuf_219 <= 0;
        FeatureBuf_220 <= 0;
        FeatureBuf_221 <= 0;
        FeatureBuf_222 <= 0;
        FeatureBuf_223 <= 0;
        FeatureBuf_224 <= 0;
        FeatureBuf_225 <= 0;
        FeatureBuf_226 <= 0;
        FeatureBuf_227 <= 0;
        FeatureBuf_228 <= 0;
        FeatureBuf_229 <= 0;
        FeatureBuf_230 <= 0;
        FeatureBuf_231 <= 0;
        FeatureBuf_232 <= 0;
        FeatureBuf_233 <= 0;
        FeatureBuf_234 <= 0;
        FeatureBuf_235 <= 0;
        FeatureBuf_236 <= 0;
        FeatureBuf_237 <= 0;
        FeatureBuf_238 <= 0;
        FeatureBuf_239 <= 0;
        FeatureBuf_240 <= 0;
        FeatureBuf_241 <= 0;
        FeatureBuf_242 <= 0;
        FeatureBuf_243 <= 0;
        FeatureBuf_244 <= 0;
        FeatureBuf_245 <= 0;
        FeatureBuf_246 <= 0;
        FeatureBuf_247 <= 0;
        FeatureBuf_248 <= 0;
        FeatureBuf_249 <= 0;
        FeatureBuf_250 <= 0;
        FeatureBuf_251 <= 0;
        FeatureBuf_252 <= 0;
        FeatureBuf_253 <= 0;
        FeatureBuf_254 <= 0;
        FeatureBuf_255 <= 0;
        FeatureBuf_256 <= 0;
        FeatureBuf_257 <= 0;
        FeatureBuf_258 <= 0;
        FeatureBuf_259 <= 0;
        FeatureBuf_260 <= 0;
        FeatureBuf_261 <= 0;
        FeatureBuf_262 <= 0;
        FeatureBuf_263 <= 0;
        FeatureBuf_264 <= 0;
        FeatureBuf_265 <= 0;
        FeatureBuf_266 <= 0;
        FeatureBuf_267 <= 0;
        FeatureBuf_268 <= 0;
        FeatureBuf_269 <= 0;
        FeatureBuf_270 <= 0;
        FeatureBuf_271 <= 0;
        FeatureBuf_272 <= 0;
        FeatureBuf_273 <= 0;
        FeatureBuf_274 <= 0;
        FeatureBuf_275 <= 0;
        FeatureBuf_276 <= 0;
        FeatureBuf_277 <= 0;
        FeatureBuf_278 <= 0;
        FeatureBuf_279 <= 0;
        FeatureBuf_280 <= 0;
        FeatureBuf_281 <= 0;
        FeatureBuf_282 <= 0;
        FeatureBuf_283 <= 0;
        FeatureBuf_284 <= 0;
        FeatureBuf_285 <= 0;
        FeatureBuf_286 <= 0;
        FeatureBuf_287 <= 0;
        FeatureBuf_288 <= 0;
        FeatureBuf_289 <= 0;
        FeatureBuf_290 <= 0;
        FeatureBuf_291 <= 0;
        FeatureBuf_292 <= 0;
        FeatureBuf_293 <= 0;
        FeatureBuf_294 <= 0;
        FeatureBuf_295 <= 0;
        FeatureBuf_296 <= 0;
        FeatureBuf_297 <= 0;
        FeatureBuf_298 <= 0;
        FeatureBuf_299 <= 0;
        FeatureBuf_300 <= 0;
        FeatureBuf_301 <= 0;
        FeatureBuf_302 <= 0;
        FeatureBuf_303 <= 0;
        FeatureBuf_304 <= 0;
        FeatureBuf_305 <= 0;
        FeatureBuf_306 <= 0;
        FeatureBuf_307 <= 0;
        FeatureBuf_308 <= 0;
        FeatureBuf_309 <= 0;
        FeatureBuf_310 <= 0;
        FeatureBuf_311 <= 0;
        FeatureBuf_312 <= 0;
        FeatureBuf_313 <= 0;
        FeatureBuf_314 <= 0;
        FeatureBuf_315 <= 0;
        FeatureBuf_316 <= 0;
        FeatureBuf_317 <= 0;
        FeatureBuf_318 <= 0;
        FeatureBuf_319 <= 0;
        FeatureBuf_320 <= 0;
        FeatureBuf_321 <= 0;
        FeatureBuf_322 <= 0;
        FeatureBuf_323 <= 0;
        FeatureBuf_324 <= 0;
        FeatureBuf_325 <= 0;
        FeatureBuf_326 <= 0;
        FeatureBuf_327 <= 0;
        FeatureBuf_328 <= 0;
        FeatureBuf_329 <= 0;
        FeatureBuf_330 <= 0;
        FeatureBuf_331 <= 0;
        FeatureBuf_332 <= 0;
        FeatureBuf_333 <= 0;
        FeatureBuf_334 <= 0;
        FeatureBuf_335 <= 0;
        FeatureBuf_336 <= 0;
        FeatureBuf_337 <= 0;
        FeatureBuf_338 <= 0;
        FeatureBuf_339 <= 0;
        FeatureBuf_340 <= 0;
        FeatureBuf_341 <= 0;
        FeatureBuf_342 <= 0;
        FeatureBuf_343 <= 0;
        FeatureBuf_344 <= 0;
        FeatureBuf_345 <= 0;
        FeatureBuf_346 <= 0;
        FeatureBuf_347 <= 0;
        FeatureBuf_348 <= 0;
        FeatureBuf_349 <= 0;
        FeatureBuf_350 <= 0;
        FeatureBuf_351 <= 0;
        FeatureBuf_352 <= 0;
        FeatureBuf_353 <= 0;
        FeatureBuf_354 <= 0;
        FeatureBuf_355 <= 0;
        FeatureBuf_356 <= 0;
        FeatureBuf_357 <= 0;
        FeatureBuf_358 <= 0;
        FeatureBuf_359 <= 0;
        FeatureBuf_360 <= 0;
        FeatureBuf_361 <= 0;
        FeatureBuf_362 <= 0;
        FeatureBuf_363 <= 0;
        FeatureBuf_364 <= 0;
        FeatureBuf_365 <= 0;
        FeatureBuf_366 <= 0;
        FeatureBuf_367 <= 0;
        FeatureBuf_368 <= 0;
        FeatureBuf_369 <= 0;
        FeatureBuf_370 <= 0;
        FeatureBuf_371 <= 0;
        FeatureBuf_372 <= 0;
        FeatureBuf_373 <= 0;
        FeatureBuf_374 <= 0;
        FeatureBuf_375 <= 0;
        FeatureBuf_376 <= 0;
        FeatureBuf_377 <= 0;
        FeatureBuf_378 <= 0;
        FeatureBuf_379 <= 0;
        FeatureBuf_380 <= 0;
        FeatureBuf_381 <= 0;
        FeatureBuf_382 <= 0;
        FeatureBuf_383 <= 0;
        FeatureBuf_384 <= 0;
        FeatureBuf_385 <= 0;
        FeatureBuf_386 <= 0;
        FeatureBuf_387 <= 0;
        FeatureBuf_388 <= 0;
        FeatureBuf_389 <= 0;
        FeatureBuf_390 <= 0;
        FeatureBuf_391 <= 0;
        FeatureBuf_392 <= 0;
        FeatureBuf_393 <= 0;
        FeatureBuf_394 <= 0;
        FeatureBuf_395 <= 0;
        FeatureBuf_396 <= 0;
        FeatureBuf_397 <= 0;
        FeatureBuf_398 <= 0;
        FeatureBuf_399 <= 0;
        FeatureBuf_400 <= 0;
        FeatureBuf_401 <= 0;
        FeatureBuf_402 <= 0;
        FeatureBuf_403 <= 0;
        FeatureBuf_404 <= 0;
        FeatureBuf_405 <= 0;
        FeatureBuf_406 <= 0;
        FeatureBuf_407 <= 0;
        FeatureBuf_408 <= 0;
        FeatureBuf_409 <= 0;
        FeatureBuf_410 <= 0;
        FeatureBuf_411 <= 0;
        FeatureBuf_412 <= 0;
        FeatureBuf_413 <= 0;
        FeatureBuf_414 <= 0;
        FeatureBuf_415 <= 0;
        FeatureBuf_416 <= 0;
        FeatureBuf_417 <= 0;
        FeatureBuf_418 <= 0;
        FeatureBuf_419 <= 0;
        FeatureBuf_420 <= 0;
        FeatureBuf_421 <= 0;
        FeatureBuf_422 <= 0;
        FeatureBuf_423 <= 0;
        FeatureBuf_424 <= 0;
        FeatureBuf_425 <= 0;
        FeatureBuf_426 <= 0;
        FeatureBuf_427 <= 0;
        FeatureBuf_428 <= 0;
        FeatureBuf_429 <= 0;
        FeatureBuf_430 <= 0;
        FeatureBuf_431 <= 0;
        FeatureBuf_432 <= 0;
        FeatureBuf_433 <= 0;
        FeatureBuf_434 <= 0;
        FeatureBuf_435 <= 0;
        FeatureBuf_436 <= 0;
        FeatureBuf_437 <= 0;
        FeatureBuf_438 <= 0;
        FeatureBuf_439 <= 0;
        FeatureBuf_440 <= 0;
        FeatureBuf_441 <= 0;
        FeatureBuf_442 <= 0;
        FeatureBuf_443 <= 0;
        FeatureBuf_444 <= 0;
        FeatureBuf_445 <= 0;
        FeatureBuf_446 <= 0;
        FeatureBuf_447 <= 0;
        FeatureBuf_448 <= 0;
        FeatureBuf_449 <= 0;
        FeatureBuf_450 <= 0;
        FeatureBuf_451 <= 0;
        FeatureBuf_452 <= 0;
        FeatureBuf_453 <= 0;
        FeatureBuf_454 <= 0;
        FeatureBuf_455 <= 0;
        FeatureBuf_456 <= 0;
        FeatureBuf_457 <= 0;
        FeatureBuf_458 <= 0;
        FeatureBuf_459 <= 0;
        FeatureBuf_460 <= 0;
        FeatureBuf_461 <= 0;
        FeatureBuf_462 <= 0;
        FeatureBuf_463 <= 0;
        FeatureBuf_464 <= 0;
        FeatureBuf_465 <= 0;
        FeatureBuf_466 <= 0;
        FeatureBuf_467 <= 0;
        FeatureBuf_468 <= 0;
        FeatureBuf_469 <= 0;
        FeatureBuf_470 <= 0;
        FeatureBuf_471 <= 0;
        FeatureBuf_472 <= 0;
        FeatureBuf_473 <= 0;
        FeatureBuf_474 <= 0;
        FeatureBuf_475 <= 0;
        FeatureBuf_476 <= 0;
        FeatureBuf_477 <= 0;
        FeatureBuf_478 <= 0;
        FeatureBuf_479 <= 0;
        FeatureBuf_480 <= 0;
        FeatureBuf_481 <= 0;
        FeatureBuf_482 <= 0;
        FeatureBuf_483 <= 0;
        FeatureBuf_484 <= 0;
        FeatureBuf_485 <= 0;
        FeatureBuf_486 <= 0;
        FeatureBuf_487 <= 0;
        FeatureBuf_488 <= 0;
        FeatureBuf_489 <= 0;
        FeatureBuf_490 <= 0;
        FeatureBuf_491 <= 0;
        FeatureBuf_492 <= 0;
        FeatureBuf_493 <= 0;
        FeatureBuf_494 <= 0;
        FeatureBuf_495 <= 0;
        FeatureBuf_496 <= 0;
        FeatureBuf_497 <= 0;
        FeatureBuf_498 <= 0;
        FeatureBuf_499 <= 0;
        FeatureBuf_500 <= 0;
        FeatureBuf_501 <= 0;
        FeatureBuf_502 <= 0;
        FeatureBuf_503 <= 0;
        FeatureBuf_504 <= 0;
        FeatureBuf_505 <= 0;
        FeatureBuf_506 <= 0;
        FeatureBuf_507 <= 0;
        FeatureBuf_508 <= 0;
        FeatureBuf_509 <= 0;
        FeatureBuf_510 <= 0;
        FeatureBuf_511 <= 0;
        FeatureBuf_512 <= 0;
        FeatureBuf_513 <= 0;
        FeatureBuf_514 <= 0;
        FeatureBuf_515 <= 0;
        FeatureBuf_516 <= 0;
        FeatureBuf_517 <= 0;
        FeatureBuf_518 <= 0;
        FeatureBuf_519 <= 0;
        FeatureBuf_520 <= 0;
        FeatureBuf_521 <= 0;
        FeatureBuf_522 <= 0;
        FeatureBuf_523 <= 0;
        FeatureBuf_524 <= 0;
        FeatureBuf_525 <= 0;
        FeatureBuf_526 <= 0;
        FeatureBuf_527 <= 0;
        FeatureBuf_528 <= 0;
        FeatureBuf_529 <= 0;
        FeatureBuf_530 <= 0;
        FeatureBuf_531 <= 0;
        FeatureBuf_532 <= 0;
        FeatureBuf_533 <= 0;
        FeatureBuf_534 <= 0;
        FeatureBuf_535 <= 0;
        FeatureBuf_536 <= 0;
        FeatureBuf_537 <= 0;
        FeatureBuf_538 <= 0;
        FeatureBuf_539 <= 0;
        FeatureBuf_540 <= 0;
        FeatureBuf_541 <= 0;
        FeatureBuf_542 <= 0;
        FeatureBuf_543 <= 0;
        FeatureBuf_544 <= 0;
        FeatureBuf_545 <= 0;
        FeatureBuf_546 <= 0;
        FeatureBuf_547 <= 0;
        FeatureBuf_548 <= 0;
        FeatureBuf_549 <= 0;
        FeatureBuf_550 <= 0;
        FeatureBuf_551 <= 0;
        FeatureBuf_552 <= 0;
        FeatureBuf_553 <= 0;
        FeatureBuf_554 <= 0;
        FeatureBuf_555 <= 0;
        FeatureBuf_556 <= 0;
        FeatureBuf_557 <= 0;
        FeatureBuf_558 <= 0;
        FeatureBuf_559 <= 0;
        FeatureBuf_560 <= 0;
        FeatureBuf_561 <= 0;
        FeatureBuf_562 <= 0;
        FeatureBuf_563 <= 0;
        FeatureBuf_564 <= 0;
        FeatureBuf_565 <= 0;
        FeatureBuf_566 <= 0;
        FeatureBuf_567 <= 0;
        FeatureBuf_568 <= 0;
        FeatureBuf_569 <= 0;
        FeatureBuf_570 <= 0;
        FeatureBuf_571 <= 0;
        FeatureBuf_572 <= 0;
        FeatureBuf_573 <= 0;
        FeatureBuf_574 <= 0;
        FeatureBuf_575 <= 0;
        FeatureBuf_576 <= 0;
        FeatureBuf_577 <= 0;
        FeatureBuf_578 <= 0;
        FeatureBuf_579 <= 0;
        FeatureBuf_580 <= 0;
        FeatureBuf_581 <= 0;
        FeatureBuf_582 <= 0;
        FeatureBuf_583 <= 0;
        FeatureBuf_584 <= 0;
        FeatureBuf_585 <= 0;
        FeatureBuf_586 <= 0;
        FeatureBuf_587 <= 0;
        FeatureBuf_588 <= 0;
        FeatureBuf_589 <= 0;
        FeatureBuf_590 <= 0;
        FeatureBuf_591 <= 0;
        FeatureBuf_592 <= 0;
        FeatureBuf_593 <= 0;
        FeatureBuf_594 <= 0;
        FeatureBuf_595 <= 0;
        FeatureBuf_596 <= 0;
        FeatureBuf_597 <= 0;
        FeatureBuf_598 <= 0;
        FeatureBuf_599 <= 0;
        FeatureBuf_600 <= 0;
        FeatureBuf_601 <= 0;
        FeatureBuf_602 <= 0;
        FeatureBuf_603 <= 0;
        FeatureBuf_604 <= 0;
        FeatureBuf_605 <= 0;
        FeatureBuf_606 <= 0;
        FeatureBuf_607 <= 0;
        FeatureBuf_608 <= 0;
        FeatureBuf_609 <= 0;
        FeatureBuf_610 <= 0;
        FeatureBuf_611 <= 0;
        FeatureBuf_612 <= 0;
        FeatureBuf_613 <= 0;
        FeatureBuf_614 <= 0;
        FeatureBuf_615 <= 0;
        FeatureBuf_616 <= 0;
        FeatureBuf_617 <= 0;
        FeatureBuf_618 <= 0;
        FeatureBuf_619 <= 0;
        FeatureBuf_620 <= 0;
        FeatureBuf_621 <= 0;
        FeatureBuf_622 <= 0;
        FeatureBuf_623 <= 0;
        FeatureBuf_624 <= 0;
        FeatureBuf_625 <= 0;
        FeatureBuf_626 <= 0;
        FeatureBuf_627 <= 0;
        FeatureBuf_628 <= 0;
        FeatureBuf_629 <= 0;
        FeatureBuf_630 <= 0;
        FeatureBuf_631 <= 0;
        FeatureBuf_632 <= 0;
        FeatureBuf_633 <= 0;
        FeatureBuf_634 <= 0;
        FeatureBuf_635 <= 0;
        FeatureBuf_636 <= 0;
        FeatureBuf_637 <= 0;
        FeatureBuf_638 <= 0;
        FeatureBuf_639 <= 0;
        FeatureBuf_640 <= 0;
        FeatureBuf_641 <= 0;
        FeatureBuf_642 <= 0;
        FeatureBuf_643 <= 0;
        FeatureBuf_644 <= 0;
        FeatureBuf_645 <= 0;
        FeatureBuf_646 <= 0;
        FeatureBuf_647 <= 0;
        FeatureBuf_648 <= 0;
        FeatureBuf_649 <= 0;
        FeatureBuf_650 <= 0;
        FeatureBuf_651 <= 0;
        FeatureBuf_652 <= 0;
        FeatureBuf_653 <= 0;
        FeatureBuf_654 <= 0;
        FeatureBuf_655 <= 0;
        FeatureBuf_656 <= 0;
        FeatureBuf_657 <= 0;
        FeatureBuf_658 <= 0;
        FeatureBuf_659 <= 0;
        FeatureBuf_660 <= 0;
        FeatureBuf_661 <= 0;
        FeatureBuf_662 <= 0;
        FeatureBuf_663 <= 0;
        FeatureBuf_664 <= 0;
        FeatureBuf_665 <= 0;
        FeatureBuf_666 <= 0;
        FeatureBuf_667 <= 0;
        FeatureBuf_668 <= 0;
        FeatureBuf_669 <= 0;
        FeatureBuf_670 <= 0;
        FeatureBuf_671 <= 0;
        FeatureBuf_672 <= 0;
        FeatureBuf_673 <= 0;
        FeatureBuf_674 <= 0;
        FeatureBuf_675 <= 0;
        FeatureBuf_676 <= 0;
        FeatureBuf_677 <= 0;
        FeatureBuf_678 <= 0;
        FeatureBuf_679 <= 0;
        FeatureBuf_680 <= 0;
        FeatureBuf_681 <= 0;
        FeatureBuf_682 <= 0;
        FeatureBuf_683 <= 0;
        FeatureBuf_684 <= 0;
        FeatureBuf_685 <= 0;
        FeatureBuf_686 <= 0;
        FeatureBuf_687 <= 0;
        FeatureBuf_688 <= 0;
        FeatureBuf_689 <= 0;
        FeatureBuf_690 <= 0;
        FeatureBuf_691 <= 0;
        FeatureBuf_692 <= 0;
        FeatureBuf_693 <= 0;
        FeatureBuf_694 <= 0;
        FeatureBuf_695 <= 0;
        FeatureBuf_696 <= 0;
        FeatureBuf_697 <= 0;
        FeatureBuf_698 <= 0;
        FeatureBuf_699 <= 0;
        FeatureBuf_700 <= 0;
        FeatureBuf_701 <= 0;
        FeatureBuf_702 <= 0;
        FeatureBuf_703 <= 0;
        FeatureBuf_704 <= 0;
        FeatureBuf_705 <= 0;
        FeatureBuf_706 <= 0;
        FeatureBuf_707 <= 0;
        FeatureBuf_708 <= 0;
        FeatureBuf_709 <= 0;
        FeatureBuf_710 <= 0;
        FeatureBuf_711 <= 0;
        FeatureBuf_712 <= 0;
        FeatureBuf_713 <= 0;
        FeatureBuf_714 <= 0;
        FeatureBuf_715 <= 0;
        FeatureBuf_716 <= 0;
        FeatureBuf_717 <= 0;
        FeatureBuf_718 <= 0;
        FeatureBuf_719 <= 0;
        FeatureBuf_720 <= 0;
        FeatureBuf_721 <= 0;
        FeatureBuf_722 <= 0;
        FeatureBuf_723 <= 0;
        FeatureBuf_724 <= 0;
        FeatureBuf_725 <= 0;
        FeatureBuf_726 <= 0;
        FeatureBuf_727 <= 0;
        FeatureBuf_728 <= 0;
        FeatureBuf_729 <= 0;
        FeatureBuf_730 <= 0;
        FeatureBuf_731 <= 0;
        FeatureBuf_732 <= 0;
        FeatureBuf_733 <= 0;
        FeatureBuf_734 <= 0;
        FeatureBuf_735 <= 0;
        FeatureBuf_736 <= 0;
        FeatureBuf_737 <= 0;
        FeatureBuf_738 <= 0;
        FeatureBuf_739 <= 0;
        FeatureBuf_740 <= 0;
        FeatureBuf_741 <= 0;
        FeatureBuf_742 <= 0;
        FeatureBuf_743 <= 0;
        FeatureBuf_744 <= 0;
        FeatureBuf_745 <= 0;
        FeatureBuf_746 <= 0;
        FeatureBuf_747 <= 0;
        FeatureBuf_748 <= 0;
        FeatureBuf_749 <= 0;
        FeatureBuf_750 <= 0;
        FeatureBuf_751 <= 0;
        FeatureBuf_752 <= 0;
        FeatureBuf_753 <= 0;
        FeatureBuf_754 <= 0;
        FeatureBuf_755 <= 0;
        FeatureBuf_756 <= 0;
        FeatureBuf_757 <= 0;
        FeatureBuf_758 <= 0;
        FeatureBuf_759 <= 0;
        FeatureBuf_760 <= 0;
        FeatureBuf_761 <= 0;
        FeatureBuf_762 <= 0;
        FeatureBuf_763 <= 0;
        FeatureBuf_764 <= 0;
        FeatureBuf_765 <= 0;
        FeatureBuf_766 <= 0;
        FeatureBuf_767 <= 0;
        FeatureBuf_768 <= 0;
        FeatureBuf_769 <= 0;
        FeatureBuf_770 <= 0;
        FeatureBuf_771 <= 0;
        FeatureBuf_772 <= 0;
        FeatureBuf_773 <= 0;
        FeatureBuf_774 <= 0;
        FeatureBuf_775 <= 0;
        FeatureBuf_776 <= 0;
        FeatureBuf_777 <= 0;
        FeatureBuf_778 <= 0;
        FeatureBuf_779 <= 0;
        FeatureBuf_780 <= 0;
        FeatureBuf_781 <= 0;
        FeatureBuf_782 <= 0;
        FeatureBuf_783 <= 0;

    end
    else if(Load) begin
        FeatureBuf_0 <= Pix_0;
        FeatureBuf_1 <= Pix_1;
        FeatureBuf_2 <= Pix_2;
        FeatureBuf_3 <= Pix_3;
        FeatureBuf_4 <= Pix_4;
        FeatureBuf_5 <= Pix_5;
        FeatureBuf_6 <= Pix_6;
        FeatureBuf_7 <= Pix_7;
        FeatureBuf_8 <= Pix_8;
        FeatureBuf_9 <= Pix_9;
        FeatureBuf_10 <= Pix_10;
        FeatureBuf_11 <= Pix_11;
        FeatureBuf_12 <= Pix_12;
        FeatureBuf_13 <= Pix_13;
        FeatureBuf_14 <= Pix_14;
        FeatureBuf_15 <= Pix_15;
        FeatureBuf_16 <= Pix_16;
        FeatureBuf_17 <= Pix_17;
        FeatureBuf_18 <= Pix_18;
        FeatureBuf_19 <= Pix_19;
        FeatureBuf_20 <= Pix_20;
        FeatureBuf_21 <= Pix_21;
        FeatureBuf_22 <= Pix_22;
        FeatureBuf_23 <= Pix_23;
        FeatureBuf_24 <= Pix_24;
        FeatureBuf_25 <= Pix_25;
        FeatureBuf_26 <= Pix_26;
        FeatureBuf_27 <= Pix_27;
        FeatureBuf_28 <= Pix_28;
        FeatureBuf_29 <= Pix_29;
        FeatureBuf_30 <= Pix_30;
        FeatureBuf_31 <= Pix_31;
        FeatureBuf_32 <= Pix_32;
        FeatureBuf_33 <= Pix_33;
        FeatureBuf_34 <= Pix_34;
        FeatureBuf_35 <= Pix_35;
        FeatureBuf_36 <= Pix_36;
        FeatureBuf_37 <= Pix_37;
        FeatureBuf_38 <= Pix_38;
        FeatureBuf_39 <= Pix_39;
        FeatureBuf_40 <= Pix_40;
        FeatureBuf_41 <= Pix_41;
        FeatureBuf_42 <= Pix_42;
        FeatureBuf_43 <= Pix_43;
        FeatureBuf_44 <= Pix_44;
        FeatureBuf_45 <= Pix_45;
        FeatureBuf_46 <= Pix_46;
        FeatureBuf_47 <= Pix_47;
        FeatureBuf_48 <= Pix_48;
        FeatureBuf_49 <= Pix_49;
        FeatureBuf_50 <= Pix_50;
        FeatureBuf_51 <= Pix_51;
        FeatureBuf_52 <= Pix_52;
        FeatureBuf_53 <= Pix_53;
        FeatureBuf_54 <= Pix_54;
        FeatureBuf_55 <= Pix_55;
        FeatureBuf_56 <= Pix_56;
        FeatureBuf_57 <= Pix_57;
        FeatureBuf_58 <= Pix_58;
        FeatureBuf_59 <= Pix_59;
        FeatureBuf_60 <= Pix_60;
        FeatureBuf_61 <= Pix_61;
        FeatureBuf_62 <= Pix_62;
        FeatureBuf_63 <= Pix_63;
        FeatureBuf_64 <= Pix_64;
        FeatureBuf_65 <= Pix_65;
        FeatureBuf_66 <= Pix_66;
        FeatureBuf_67 <= Pix_67;
        FeatureBuf_68 <= Pix_68;
        FeatureBuf_69 <= Pix_69;
        FeatureBuf_70 <= Pix_70;
        FeatureBuf_71 <= Pix_71;
        FeatureBuf_72 <= Pix_72;
        FeatureBuf_73 <= Pix_73;
        FeatureBuf_74 <= Pix_74;
        FeatureBuf_75 <= Pix_75;
        FeatureBuf_76 <= Pix_76;
        FeatureBuf_77 <= Pix_77;
        FeatureBuf_78 <= Pix_78;
        FeatureBuf_79 <= Pix_79;
        FeatureBuf_80 <= Pix_80;
        FeatureBuf_81 <= Pix_81;
        FeatureBuf_82 <= Pix_82;
        FeatureBuf_83 <= Pix_83;
        FeatureBuf_84 <= Pix_84;
        FeatureBuf_85 <= Pix_85;
        FeatureBuf_86 <= Pix_86;
        FeatureBuf_87 <= Pix_87;
        FeatureBuf_88 <= Pix_88;
        FeatureBuf_89 <= Pix_89;
        FeatureBuf_90 <= Pix_90;
        FeatureBuf_91 <= Pix_91;
        FeatureBuf_92 <= Pix_92;
        FeatureBuf_93 <= Pix_93;
        FeatureBuf_94 <= Pix_94;
        FeatureBuf_95 <= Pix_95;
        FeatureBuf_96 <= Pix_96;
        FeatureBuf_97 <= Pix_97;
        FeatureBuf_98 <= Pix_98;
        FeatureBuf_99 <= Pix_99;
        FeatureBuf_100 <= Pix_100;
        FeatureBuf_101 <= Pix_101;
        FeatureBuf_102 <= Pix_102;
        FeatureBuf_103 <= Pix_103;
        FeatureBuf_104 <= Pix_104;
        FeatureBuf_105 <= Pix_105;
        FeatureBuf_106 <= Pix_106;
        FeatureBuf_107 <= Pix_107;
        FeatureBuf_108 <= Pix_108;
        FeatureBuf_109 <= Pix_109;
        FeatureBuf_110 <= Pix_110;
        FeatureBuf_111 <= Pix_111;
        FeatureBuf_112 <= Pix_112;
        FeatureBuf_113 <= Pix_113;
        FeatureBuf_114 <= Pix_114;
        FeatureBuf_115 <= Pix_115;
        FeatureBuf_116 <= Pix_116;
        FeatureBuf_117 <= Pix_117;
        FeatureBuf_118 <= Pix_118;
        FeatureBuf_119 <= Pix_119;
        FeatureBuf_120 <= Pix_120;
        FeatureBuf_121 <= Pix_121;
        FeatureBuf_122 <= Pix_122;
        FeatureBuf_123 <= Pix_123;
        FeatureBuf_124 <= Pix_124;
        FeatureBuf_125 <= Pix_125;
        FeatureBuf_126 <= Pix_126;
        FeatureBuf_127 <= Pix_127;
        FeatureBuf_128 <= Pix_128;
        FeatureBuf_129 <= Pix_129;
        FeatureBuf_130 <= Pix_130;
        FeatureBuf_131 <= Pix_131;
        FeatureBuf_132 <= Pix_132;
        FeatureBuf_133 <= Pix_133;
        FeatureBuf_134 <= Pix_134;
        FeatureBuf_135 <= Pix_135;
        FeatureBuf_136 <= Pix_136;
        FeatureBuf_137 <= Pix_137;
        FeatureBuf_138 <= Pix_138;
        FeatureBuf_139 <= Pix_139;
        FeatureBuf_140 <= Pix_140;
        FeatureBuf_141 <= Pix_141;
        FeatureBuf_142 <= Pix_142;
        FeatureBuf_143 <= Pix_143;
        FeatureBuf_144 <= Pix_144;
        FeatureBuf_145 <= Pix_145;
        FeatureBuf_146 <= Pix_146;
        FeatureBuf_147 <= Pix_147;
        FeatureBuf_148 <= Pix_148;
        FeatureBuf_149 <= Pix_149;
        FeatureBuf_150 <= Pix_150;
        FeatureBuf_151 <= Pix_151;
        FeatureBuf_152 <= Pix_152;
        FeatureBuf_153 <= Pix_153;
        FeatureBuf_154 <= Pix_154;
        FeatureBuf_155 <= Pix_155;
        FeatureBuf_156 <= Pix_156;
        FeatureBuf_157 <= Pix_157;
        FeatureBuf_158 <= Pix_158;
        FeatureBuf_159 <= Pix_159;
        FeatureBuf_160 <= Pix_160;
        FeatureBuf_161 <= Pix_161;
        FeatureBuf_162 <= Pix_162;
        FeatureBuf_163 <= Pix_163;
        FeatureBuf_164 <= Pix_164;
        FeatureBuf_165 <= Pix_165;
        FeatureBuf_166 <= Pix_166;
        FeatureBuf_167 <= Pix_167;
        FeatureBuf_168 <= Pix_168;
        FeatureBuf_169 <= Pix_169;
        FeatureBuf_170 <= Pix_170;
        FeatureBuf_171 <= Pix_171;
        FeatureBuf_172 <= Pix_172;
        FeatureBuf_173 <= Pix_173;
        FeatureBuf_174 <= Pix_174;
        FeatureBuf_175 <= Pix_175;
        FeatureBuf_176 <= Pix_176;
        FeatureBuf_177 <= Pix_177;
        FeatureBuf_178 <= Pix_178;
        FeatureBuf_179 <= Pix_179;
        FeatureBuf_180 <= Pix_180;
        FeatureBuf_181 <= Pix_181;
        FeatureBuf_182 <= Pix_182;
        FeatureBuf_183 <= Pix_183;
        FeatureBuf_184 <= Pix_184;
        FeatureBuf_185 <= Pix_185;
        FeatureBuf_186 <= Pix_186;
        FeatureBuf_187 <= Pix_187;
        FeatureBuf_188 <= Pix_188;
        FeatureBuf_189 <= Pix_189;
        FeatureBuf_190 <= Pix_190;
        FeatureBuf_191 <= Pix_191;
        FeatureBuf_192 <= Pix_192;
        FeatureBuf_193 <= Pix_193;
        FeatureBuf_194 <= Pix_194;
        FeatureBuf_195 <= Pix_195;
        FeatureBuf_196 <= Pix_196;
        FeatureBuf_197 <= Pix_197;
        FeatureBuf_198 <= Pix_198;
        FeatureBuf_199 <= Pix_199;
        FeatureBuf_200 <= Pix_200;
        FeatureBuf_201 <= Pix_201;
        FeatureBuf_202 <= Pix_202;
        FeatureBuf_203 <= Pix_203;
        FeatureBuf_204 <= Pix_204;
        FeatureBuf_205 <= Pix_205;
        FeatureBuf_206 <= Pix_206;
        FeatureBuf_207 <= Pix_207;
        FeatureBuf_208 <= Pix_208;
        FeatureBuf_209 <= Pix_209;
        FeatureBuf_210 <= Pix_210;
        FeatureBuf_211 <= Pix_211;
        FeatureBuf_212 <= Pix_212;
        FeatureBuf_213 <= Pix_213;
        FeatureBuf_214 <= Pix_214;
        FeatureBuf_215 <= Pix_215;
        FeatureBuf_216 <= Pix_216;
        FeatureBuf_217 <= Pix_217;
        FeatureBuf_218 <= Pix_218;
        FeatureBuf_219 <= Pix_219;
        FeatureBuf_220 <= Pix_220;
        FeatureBuf_221 <= Pix_221;
        FeatureBuf_222 <= Pix_222;
        FeatureBuf_223 <= Pix_223;
        FeatureBuf_224 <= Pix_224;
        FeatureBuf_225 <= Pix_225;
        FeatureBuf_226 <= Pix_226;
        FeatureBuf_227 <= Pix_227;
        FeatureBuf_228 <= Pix_228;
        FeatureBuf_229 <= Pix_229;
        FeatureBuf_230 <= Pix_230;
        FeatureBuf_231 <= Pix_231;
        FeatureBuf_232 <= Pix_232;
        FeatureBuf_233 <= Pix_233;
        FeatureBuf_234 <= Pix_234;
        FeatureBuf_235 <= Pix_235;
        FeatureBuf_236 <= Pix_236;
        FeatureBuf_237 <= Pix_237;
        FeatureBuf_238 <= Pix_238;
        FeatureBuf_239 <= Pix_239;
        FeatureBuf_240 <= Pix_240;
        FeatureBuf_241 <= Pix_241;
        FeatureBuf_242 <= Pix_242;
        FeatureBuf_243 <= Pix_243;
        FeatureBuf_244 <= Pix_244;
        FeatureBuf_245 <= Pix_245;
        FeatureBuf_246 <= Pix_246;
        FeatureBuf_247 <= Pix_247;
        FeatureBuf_248 <= Pix_248;
        FeatureBuf_249 <= Pix_249;
        FeatureBuf_250 <= Pix_250;
        FeatureBuf_251 <= Pix_251;
        FeatureBuf_252 <= Pix_252;
        FeatureBuf_253 <= Pix_253;
        FeatureBuf_254 <= Pix_254;
        FeatureBuf_255 <= Pix_255;
        FeatureBuf_256 <= Pix_256;
        FeatureBuf_257 <= Pix_257;
        FeatureBuf_258 <= Pix_258;
        FeatureBuf_259 <= Pix_259;
        FeatureBuf_260 <= Pix_260;
        FeatureBuf_261 <= Pix_261;
        FeatureBuf_262 <= Pix_262;
        FeatureBuf_263 <= Pix_263;
        FeatureBuf_264 <= Pix_264;
        FeatureBuf_265 <= Pix_265;
        FeatureBuf_266 <= Pix_266;
        FeatureBuf_267 <= Pix_267;
        FeatureBuf_268 <= Pix_268;
        FeatureBuf_269 <= Pix_269;
        FeatureBuf_270 <= Pix_270;
        FeatureBuf_271 <= Pix_271;
        FeatureBuf_272 <= Pix_272;
        FeatureBuf_273 <= Pix_273;
        FeatureBuf_274 <= Pix_274;
        FeatureBuf_275 <= Pix_275;
        FeatureBuf_276 <= Pix_276;
        FeatureBuf_277 <= Pix_277;
        FeatureBuf_278 <= Pix_278;
        FeatureBuf_279 <= Pix_279;
        FeatureBuf_280 <= Pix_280;
        FeatureBuf_281 <= Pix_281;
        FeatureBuf_282 <= Pix_282;
        FeatureBuf_283 <= Pix_283;
        FeatureBuf_284 <= Pix_284;
        FeatureBuf_285 <= Pix_285;
        FeatureBuf_286 <= Pix_286;
        FeatureBuf_287 <= Pix_287;
        FeatureBuf_288 <= Pix_288;
        FeatureBuf_289 <= Pix_289;
        FeatureBuf_290 <= Pix_290;
        FeatureBuf_291 <= Pix_291;
        FeatureBuf_292 <= Pix_292;
        FeatureBuf_293 <= Pix_293;
        FeatureBuf_294 <= Pix_294;
        FeatureBuf_295 <= Pix_295;
        FeatureBuf_296 <= Pix_296;
        FeatureBuf_297 <= Pix_297;
        FeatureBuf_298 <= Pix_298;
        FeatureBuf_299 <= Pix_299;
        FeatureBuf_300 <= Pix_300;
        FeatureBuf_301 <= Pix_301;
        FeatureBuf_302 <= Pix_302;
        FeatureBuf_303 <= Pix_303;
        FeatureBuf_304 <= Pix_304;
        FeatureBuf_305 <= Pix_305;
        FeatureBuf_306 <= Pix_306;
        FeatureBuf_307 <= Pix_307;
        FeatureBuf_308 <= Pix_308;
        FeatureBuf_309 <= Pix_309;
        FeatureBuf_310 <= Pix_310;
        FeatureBuf_311 <= Pix_311;
        FeatureBuf_312 <= Pix_312;
        FeatureBuf_313 <= Pix_313;
        FeatureBuf_314 <= Pix_314;
        FeatureBuf_315 <= Pix_315;
        FeatureBuf_316 <= Pix_316;
        FeatureBuf_317 <= Pix_317;
        FeatureBuf_318 <= Pix_318;
        FeatureBuf_319 <= Pix_319;
        FeatureBuf_320 <= Pix_320;
        FeatureBuf_321 <= Pix_321;
        FeatureBuf_322 <= Pix_322;
        FeatureBuf_323 <= Pix_323;
        FeatureBuf_324 <= Pix_324;
        FeatureBuf_325 <= Pix_325;
        FeatureBuf_326 <= Pix_326;
        FeatureBuf_327 <= Pix_327;
        FeatureBuf_328 <= Pix_328;
        FeatureBuf_329 <= Pix_329;
        FeatureBuf_330 <= Pix_330;
        FeatureBuf_331 <= Pix_331;
        FeatureBuf_332 <= Pix_332;
        FeatureBuf_333 <= Pix_333;
        FeatureBuf_334 <= Pix_334;
        FeatureBuf_335 <= Pix_335;
        FeatureBuf_336 <= Pix_336;
        FeatureBuf_337 <= Pix_337;
        FeatureBuf_338 <= Pix_338;
        FeatureBuf_339 <= Pix_339;
        FeatureBuf_340 <= Pix_340;
        FeatureBuf_341 <= Pix_341;
        FeatureBuf_342 <= Pix_342;
        FeatureBuf_343 <= Pix_343;
        FeatureBuf_344 <= Pix_344;
        FeatureBuf_345 <= Pix_345;
        FeatureBuf_346 <= Pix_346;
        FeatureBuf_347 <= Pix_347;
        FeatureBuf_348 <= Pix_348;
        FeatureBuf_349 <= Pix_349;
        FeatureBuf_350 <= Pix_350;
        FeatureBuf_351 <= Pix_351;
        FeatureBuf_352 <= Pix_352;
        FeatureBuf_353 <= Pix_353;
        FeatureBuf_354 <= Pix_354;
        FeatureBuf_355 <= Pix_355;
        FeatureBuf_356 <= Pix_356;
        FeatureBuf_357 <= Pix_357;
        FeatureBuf_358 <= Pix_358;
        FeatureBuf_359 <= Pix_359;
        FeatureBuf_360 <= Pix_360;
        FeatureBuf_361 <= Pix_361;
        FeatureBuf_362 <= Pix_362;
        FeatureBuf_363 <= Pix_363;
        FeatureBuf_364 <= Pix_364;
        FeatureBuf_365 <= Pix_365;
        FeatureBuf_366 <= Pix_366;
        FeatureBuf_367 <= Pix_367;
        FeatureBuf_368 <= Pix_368;
        FeatureBuf_369 <= Pix_369;
        FeatureBuf_370 <= Pix_370;
        FeatureBuf_371 <= Pix_371;
        FeatureBuf_372 <= Pix_372;
        FeatureBuf_373 <= Pix_373;
        FeatureBuf_374 <= Pix_374;
        FeatureBuf_375 <= Pix_375;
        FeatureBuf_376 <= Pix_376;
        FeatureBuf_377 <= Pix_377;
        FeatureBuf_378 <= Pix_378;
        FeatureBuf_379 <= Pix_379;
        FeatureBuf_380 <= Pix_380;
        FeatureBuf_381 <= Pix_381;
        FeatureBuf_382 <= Pix_382;
        FeatureBuf_383 <= Pix_383;
        FeatureBuf_384 <= Pix_384;
        FeatureBuf_385 <= Pix_385;
        FeatureBuf_386 <= Pix_386;
        FeatureBuf_387 <= Pix_387;
        FeatureBuf_388 <= Pix_388;
        FeatureBuf_389 <= Pix_389;
        FeatureBuf_390 <= Pix_390;
        FeatureBuf_391 <= Pix_391;
        FeatureBuf_392 <= Pix_392;
        FeatureBuf_393 <= Pix_393;
        FeatureBuf_394 <= Pix_394;
        FeatureBuf_395 <= Pix_395;
        FeatureBuf_396 <= Pix_396;
        FeatureBuf_397 <= Pix_397;
        FeatureBuf_398 <= Pix_398;
        FeatureBuf_399 <= Pix_399;
        FeatureBuf_400 <= Pix_400;
        FeatureBuf_401 <= Pix_401;
        FeatureBuf_402 <= Pix_402;
        FeatureBuf_403 <= Pix_403;
        FeatureBuf_404 <= Pix_404;
        FeatureBuf_405 <= Pix_405;
        FeatureBuf_406 <= Pix_406;
        FeatureBuf_407 <= Pix_407;
        FeatureBuf_408 <= Pix_408;
        FeatureBuf_409 <= Pix_409;
        FeatureBuf_410 <= Pix_410;
        FeatureBuf_411 <= Pix_411;
        FeatureBuf_412 <= Pix_412;
        FeatureBuf_413 <= Pix_413;
        FeatureBuf_414 <= Pix_414;
        FeatureBuf_415 <= Pix_415;
        FeatureBuf_416 <= Pix_416;
        FeatureBuf_417 <= Pix_417;
        FeatureBuf_418 <= Pix_418;
        FeatureBuf_419 <= Pix_419;
        FeatureBuf_420 <= Pix_420;
        FeatureBuf_421 <= Pix_421;
        FeatureBuf_422 <= Pix_422;
        FeatureBuf_423 <= Pix_423;
        FeatureBuf_424 <= Pix_424;
        FeatureBuf_425 <= Pix_425;
        FeatureBuf_426 <= Pix_426;
        FeatureBuf_427 <= Pix_427;
        FeatureBuf_428 <= Pix_428;
        FeatureBuf_429 <= Pix_429;
        FeatureBuf_430 <= Pix_430;
        FeatureBuf_431 <= Pix_431;
        FeatureBuf_432 <= Pix_432;
        FeatureBuf_433 <= Pix_433;
        FeatureBuf_434 <= Pix_434;
        FeatureBuf_435 <= Pix_435;
        FeatureBuf_436 <= Pix_436;
        FeatureBuf_437 <= Pix_437;
        FeatureBuf_438 <= Pix_438;
        FeatureBuf_439 <= Pix_439;
        FeatureBuf_440 <= Pix_440;
        FeatureBuf_441 <= Pix_441;
        FeatureBuf_442 <= Pix_442;
        FeatureBuf_443 <= Pix_443;
        FeatureBuf_444 <= Pix_444;
        FeatureBuf_445 <= Pix_445;
        FeatureBuf_446 <= Pix_446;
        FeatureBuf_447 <= Pix_447;
        FeatureBuf_448 <= Pix_448;
        FeatureBuf_449 <= Pix_449;
        FeatureBuf_450 <= Pix_450;
        FeatureBuf_451 <= Pix_451;
        FeatureBuf_452 <= Pix_452;
        FeatureBuf_453 <= Pix_453;
        FeatureBuf_454 <= Pix_454;
        FeatureBuf_455 <= Pix_455;
        FeatureBuf_456 <= Pix_456;
        FeatureBuf_457 <= Pix_457;
        FeatureBuf_458 <= Pix_458;
        FeatureBuf_459 <= Pix_459;
        FeatureBuf_460 <= Pix_460;
        FeatureBuf_461 <= Pix_461;
        FeatureBuf_462 <= Pix_462;
        FeatureBuf_463 <= Pix_463;
        FeatureBuf_464 <= Pix_464;
        FeatureBuf_465 <= Pix_465;
        FeatureBuf_466 <= Pix_466;
        FeatureBuf_467 <= Pix_467;
        FeatureBuf_468 <= Pix_468;
        FeatureBuf_469 <= Pix_469;
        FeatureBuf_470 <= Pix_470;
        FeatureBuf_471 <= Pix_471;
        FeatureBuf_472 <= Pix_472;
        FeatureBuf_473 <= Pix_473;
        FeatureBuf_474 <= Pix_474;
        FeatureBuf_475 <= Pix_475;
        FeatureBuf_476 <= Pix_476;
        FeatureBuf_477 <= Pix_477;
        FeatureBuf_478 <= Pix_478;
        FeatureBuf_479 <= Pix_479;
        FeatureBuf_480 <= Pix_480;
        FeatureBuf_481 <= Pix_481;
        FeatureBuf_482 <= Pix_482;
        FeatureBuf_483 <= Pix_483;
        FeatureBuf_484 <= Pix_484;
        FeatureBuf_485 <= Pix_485;
        FeatureBuf_486 <= Pix_486;
        FeatureBuf_487 <= Pix_487;
        FeatureBuf_488 <= Pix_488;
        FeatureBuf_489 <= Pix_489;
        FeatureBuf_490 <= Pix_490;
        FeatureBuf_491 <= Pix_491;
        FeatureBuf_492 <= Pix_492;
        FeatureBuf_493 <= Pix_493;
        FeatureBuf_494 <= Pix_494;
        FeatureBuf_495 <= Pix_495;
        FeatureBuf_496 <= Pix_496;
        FeatureBuf_497 <= Pix_497;
        FeatureBuf_498 <= Pix_498;
        FeatureBuf_499 <= Pix_499;
        FeatureBuf_500 <= Pix_500;
        FeatureBuf_501 <= Pix_501;
        FeatureBuf_502 <= Pix_502;
        FeatureBuf_503 <= Pix_503;
        FeatureBuf_504 <= Pix_504;
        FeatureBuf_505 <= Pix_505;
        FeatureBuf_506 <= Pix_506;
        FeatureBuf_507 <= Pix_507;
        FeatureBuf_508 <= Pix_508;
        FeatureBuf_509 <= Pix_509;
        FeatureBuf_510 <= Pix_510;
        FeatureBuf_511 <= Pix_511;
        FeatureBuf_512 <= Pix_512;
        FeatureBuf_513 <= Pix_513;
        FeatureBuf_514 <= Pix_514;
        FeatureBuf_515 <= Pix_515;
        FeatureBuf_516 <= Pix_516;
        FeatureBuf_517 <= Pix_517;
        FeatureBuf_518 <= Pix_518;
        FeatureBuf_519 <= Pix_519;
        FeatureBuf_520 <= Pix_520;
        FeatureBuf_521 <= Pix_521;
        FeatureBuf_522 <= Pix_522;
        FeatureBuf_523 <= Pix_523;
        FeatureBuf_524 <= Pix_524;
        FeatureBuf_525 <= Pix_525;
        FeatureBuf_526 <= Pix_526;
        FeatureBuf_527 <= Pix_527;
        FeatureBuf_528 <= Pix_528;
        FeatureBuf_529 <= Pix_529;
        FeatureBuf_530 <= Pix_530;
        FeatureBuf_531 <= Pix_531;
        FeatureBuf_532 <= Pix_532;
        FeatureBuf_533 <= Pix_533;
        FeatureBuf_534 <= Pix_534;
        FeatureBuf_535 <= Pix_535;
        FeatureBuf_536 <= Pix_536;
        FeatureBuf_537 <= Pix_537;
        FeatureBuf_538 <= Pix_538;
        FeatureBuf_539 <= Pix_539;
        FeatureBuf_540 <= Pix_540;
        FeatureBuf_541 <= Pix_541;
        FeatureBuf_542 <= Pix_542;
        FeatureBuf_543 <= Pix_543;
        FeatureBuf_544 <= Pix_544;
        FeatureBuf_545 <= Pix_545;
        FeatureBuf_546 <= Pix_546;
        FeatureBuf_547 <= Pix_547;
        FeatureBuf_548 <= Pix_548;
        FeatureBuf_549 <= Pix_549;
        FeatureBuf_550 <= Pix_550;
        FeatureBuf_551 <= Pix_551;
        FeatureBuf_552 <= Pix_552;
        FeatureBuf_553 <= Pix_553;
        FeatureBuf_554 <= Pix_554;
        FeatureBuf_555 <= Pix_555;
        FeatureBuf_556 <= Pix_556;
        FeatureBuf_557 <= Pix_557;
        FeatureBuf_558 <= Pix_558;
        FeatureBuf_559 <= Pix_559;
        FeatureBuf_560 <= Pix_560;
        FeatureBuf_561 <= Pix_561;
        FeatureBuf_562 <= Pix_562;
        FeatureBuf_563 <= Pix_563;
        FeatureBuf_564 <= Pix_564;
        FeatureBuf_565 <= Pix_565;
        FeatureBuf_566 <= Pix_566;
        FeatureBuf_567 <= Pix_567;
        FeatureBuf_568 <= Pix_568;
        FeatureBuf_569 <= Pix_569;
        FeatureBuf_570 <= Pix_570;
        FeatureBuf_571 <= Pix_571;
        FeatureBuf_572 <= Pix_572;
        FeatureBuf_573 <= Pix_573;
        FeatureBuf_574 <= Pix_574;
        FeatureBuf_575 <= Pix_575;
        FeatureBuf_576 <= Pix_576;
        FeatureBuf_577 <= Pix_577;
        FeatureBuf_578 <= Pix_578;
        FeatureBuf_579 <= Pix_579;
        FeatureBuf_580 <= Pix_580;
        FeatureBuf_581 <= Pix_581;
        FeatureBuf_582 <= Pix_582;
        FeatureBuf_583 <= Pix_583;
        FeatureBuf_584 <= Pix_584;
        FeatureBuf_585 <= Pix_585;
        FeatureBuf_586 <= Pix_586;
        FeatureBuf_587 <= Pix_587;
        FeatureBuf_588 <= Pix_588;
        FeatureBuf_589 <= Pix_589;
        FeatureBuf_590 <= Pix_590;
        FeatureBuf_591 <= Pix_591;
        FeatureBuf_592 <= Pix_592;
        FeatureBuf_593 <= Pix_593;
        FeatureBuf_594 <= Pix_594;
        FeatureBuf_595 <= Pix_595;
        FeatureBuf_596 <= Pix_596;
        FeatureBuf_597 <= Pix_597;
        FeatureBuf_598 <= Pix_598;
        FeatureBuf_599 <= Pix_599;
        FeatureBuf_600 <= Pix_600;
        FeatureBuf_601 <= Pix_601;
        FeatureBuf_602 <= Pix_602;
        FeatureBuf_603 <= Pix_603;
        FeatureBuf_604 <= Pix_604;
        FeatureBuf_605 <= Pix_605;
        FeatureBuf_606 <= Pix_606;
        FeatureBuf_607 <= Pix_607;
        FeatureBuf_608 <= Pix_608;
        FeatureBuf_609 <= Pix_609;
        FeatureBuf_610 <= Pix_610;
        FeatureBuf_611 <= Pix_611;
        FeatureBuf_612 <= Pix_612;
        FeatureBuf_613 <= Pix_613;
        FeatureBuf_614 <= Pix_614;
        FeatureBuf_615 <= Pix_615;
        FeatureBuf_616 <= Pix_616;
        FeatureBuf_617 <= Pix_617;
        FeatureBuf_618 <= Pix_618;
        FeatureBuf_619 <= Pix_619;
        FeatureBuf_620 <= Pix_620;
        FeatureBuf_621 <= Pix_621;
        FeatureBuf_622 <= Pix_622;
        FeatureBuf_623 <= Pix_623;
        FeatureBuf_624 <= Pix_624;
        FeatureBuf_625 <= Pix_625;
        FeatureBuf_626 <= Pix_626;
        FeatureBuf_627 <= Pix_627;
        FeatureBuf_628 <= Pix_628;
        FeatureBuf_629 <= Pix_629;
        FeatureBuf_630 <= Pix_630;
        FeatureBuf_631 <= Pix_631;
        FeatureBuf_632 <= Pix_632;
        FeatureBuf_633 <= Pix_633;
        FeatureBuf_634 <= Pix_634;
        FeatureBuf_635 <= Pix_635;
        FeatureBuf_636 <= Pix_636;
        FeatureBuf_637 <= Pix_637;
        FeatureBuf_638 <= Pix_638;
        FeatureBuf_639 <= Pix_639;
        FeatureBuf_640 <= Pix_640;
        FeatureBuf_641 <= Pix_641;
        FeatureBuf_642 <= Pix_642;
        FeatureBuf_643 <= Pix_643;
        FeatureBuf_644 <= Pix_644;
        FeatureBuf_645 <= Pix_645;
        FeatureBuf_646 <= Pix_646;
        FeatureBuf_647 <= Pix_647;
        FeatureBuf_648 <= Pix_648;
        FeatureBuf_649 <= Pix_649;
        FeatureBuf_650 <= Pix_650;
        FeatureBuf_651 <= Pix_651;
        FeatureBuf_652 <= Pix_652;
        FeatureBuf_653 <= Pix_653;
        FeatureBuf_654 <= Pix_654;
        FeatureBuf_655 <= Pix_655;
        FeatureBuf_656 <= Pix_656;
        FeatureBuf_657 <= Pix_657;
        FeatureBuf_658 <= Pix_658;
        FeatureBuf_659 <= Pix_659;
        FeatureBuf_660 <= Pix_660;
        FeatureBuf_661 <= Pix_661;
        FeatureBuf_662 <= Pix_662;
        FeatureBuf_663 <= Pix_663;
        FeatureBuf_664 <= Pix_664;
        FeatureBuf_665 <= Pix_665;
        FeatureBuf_666 <= Pix_666;
        FeatureBuf_667 <= Pix_667;
        FeatureBuf_668 <= Pix_668;
        FeatureBuf_669 <= Pix_669;
        FeatureBuf_670 <= Pix_670;
        FeatureBuf_671 <= Pix_671;
        FeatureBuf_672 <= Pix_672;
        FeatureBuf_673 <= Pix_673;
        FeatureBuf_674 <= Pix_674;
        FeatureBuf_675 <= Pix_675;
        FeatureBuf_676 <= Pix_676;
        FeatureBuf_677 <= Pix_677;
        FeatureBuf_678 <= Pix_678;
        FeatureBuf_679 <= Pix_679;
        FeatureBuf_680 <= Pix_680;
        FeatureBuf_681 <= Pix_681;
        FeatureBuf_682 <= Pix_682;
        FeatureBuf_683 <= Pix_683;
        FeatureBuf_684 <= Pix_684;
        FeatureBuf_685 <= Pix_685;
        FeatureBuf_686 <= Pix_686;
        FeatureBuf_687 <= Pix_687;
        FeatureBuf_688 <= Pix_688;
        FeatureBuf_689 <= Pix_689;
        FeatureBuf_690 <= Pix_690;
        FeatureBuf_691 <= Pix_691;
        FeatureBuf_692 <= Pix_692;
        FeatureBuf_693 <= Pix_693;
        FeatureBuf_694 <= Pix_694;
        FeatureBuf_695 <= Pix_695;
        FeatureBuf_696 <= Pix_696;
        FeatureBuf_697 <= Pix_697;
        FeatureBuf_698 <= Pix_698;
        FeatureBuf_699 <= Pix_699;
        FeatureBuf_700 <= Pix_700;
        FeatureBuf_701 <= Pix_701;
        FeatureBuf_702 <= Pix_702;
        FeatureBuf_703 <= Pix_703;
        FeatureBuf_704 <= Pix_704;
        FeatureBuf_705 <= Pix_705;
        FeatureBuf_706 <= Pix_706;
        FeatureBuf_707 <= Pix_707;
        FeatureBuf_708 <= Pix_708;
        FeatureBuf_709 <= Pix_709;
        FeatureBuf_710 <= Pix_710;
        FeatureBuf_711 <= Pix_711;
        FeatureBuf_712 <= Pix_712;
        FeatureBuf_713 <= Pix_713;
        FeatureBuf_714 <= Pix_714;
        FeatureBuf_715 <= Pix_715;
        FeatureBuf_716 <= Pix_716;
        FeatureBuf_717 <= Pix_717;
        FeatureBuf_718 <= Pix_718;
        FeatureBuf_719 <= Pix_719;
        FeatureBuf_720 <= Pix_720;
        FeatureBuf_721 <= Pix_721;
        FeatureBuf_722 <= Pix_722;
        FeatureBuf_723 <= Pix_723;
        FeatureBuf_724 <= Pix_724;
        FeatureBuf_725 <= Pix_725;
        FeatureBuf_726 <= Pix_726;
        FeatureBuf_727 <= Pix_727;
        FeatureBuf_728 <= Pix_728;
        FeatureBuf_729 <= Pix_729;
        FeatureBuf_730 <= Pix_730;
        FeatureBuf_731 <= Pix_731;
        FeatureBuf_732 <= Pix_732;
        FeatureBuf_733 <= Pix_733;
        FeatureBuf_734 <= Pix_734;
        FeatureBuf_735 <= Pix_735;
        FeatureBuf_736 <= Pix_736;
        FeatureBuf_737 <= Pix_737;
        FeatureBuf_738 <= Pix_738;
        FeatureBuf_739 <= Pix_739;
        FeatureBuf_740 <= Pix_740;
        FeatureBuf_741 <= Pix_741;
        FeatureBuf_742 <= Pix_742;
        FeatureBuf_743 <= Pix_743;
        FeatureBuf_744 <= Pix_744;
        FeatureBuf_745 <= Pix_745;
        FeatureBuf_746 <= Pix_746;
        FeatureBuf_747 <= Pix_747;
        FeatureBuf_748 <= Pix_748;
        FeatureBuf_749 <= Pix_749;
        FeatureBuf_750 <= Pix_750;
        FeatureBuf_751 <= Pix_751;
        FeatureBuf_752 <= Pix_752;
        FeatureBuf_753 <= Pix_753;
        FeatureBuf_754 <= Pix_754;
        FeatureBuf_755 <= Pix_755;
        FeatureBuf_756 <= Pix_756;
        FeatureBuf_757 <= Pix_757;
        FeatureBuf_758 <= Pix_758;
        FeatureBuf_759 <= Pix_759;
        FeatureBuf_760 <= Pix_760;
        FeatureBuf_761 <= Pix_761;
        FeatureBuf_762 <= Pix_762;
        FeatureBuf_763 <= Pix_763;
        FeatureBuf_764 <= Pix_764;
        FeatureBuf_765 <= Pix_765;
        FeatureBuf_766 <= Pix_766;
        FeatureBuf_767 <= Pix_767;
        FeatureBuf_768 <= Pix_768;
        FeatureBuf_769 <= Pix_769;
        FeatureBuf_770 <= Pix_770;
        FeatureBuf_771 <= Pix_771;
        FeatureBuf_772 <= Pix_772;
        FeatureBuf_773 <= Pix_773;
        FeatureBuf_774 <= Pix_774;
        FeatureBuf_775 <= Pix_775;
        FeatureBuf_776 <= Pix_776;
        FeatureBuf_777 <= Pix_777;
        FeatureBuf_778 <= Pix_778;
        FeatureBuf_779 <= Pix_779;
        FeatureBuf_780 <= Pix_780;
        FeatureBuf_781 <= Pix_781;
        FeatureBuf_782 <= Pix_782;
        FeatureBuf_783 <= Pix_783;


    end
end

always@(posedge clk, negedge GlobalReset)begin
    if(!GlobalReset)begin
        Res0 <= 0;
        Res1 <= 0;
        Res2 <= 0;
        Res3 <= 0;
        Res4 <= 0;
        Res5 <= 0;
        Res6 <= 0;
        Res7 <= 0;
        Res8 <= 0;
        Res9 <= 0;
    end
    else begin
        Res0 <= Res0_n;
        Res1 <= Res1_n;
        Res2 <= Res2_n;
        Res3 <= Res3_n;
        Res4 <= Res4_n;
        Res5 <= Res5_n;
        Res6 <= Res6_n;
        Res7 <= Res7_n;
        Res8 <= Res8_n;
        Res9 <= Res9_n;
    end
end

always@(posedge clk, negedge GlobalReset)begin
    if(!GlobalReset)begin
        Res_0_0 <= 0;
        Res_0_1 <= 0;
        Res_0_2 <= 0;
        Res_0_3 <= 0;
        Res_0_4 <= 0;
        Res_0_5 <= 0;
        Res_0_6 <= 0;
        Res_0_7 <= 0;
        Res_1_0 <= 0;
        Res_1_1 <= 0;
        Res_1_2 <= 0;
        Res_1_3 <= 0;
        Res_1_4 <= 0;
        Res_1_5 <= 0;
        Res_1_6 <= 0;
        Res_1_7 <= 0;
        Res_2_0 <= 0;
        Res_2_1 <= 0;
        Res_2_2 <= 0;
        Res_2_3 <= 0;
        Res_2_4 <= 0;
        Res_2_5 <= 0;
        Res_2_6 <= 0;
        Res_2_7 <= 0;
        Res_3_0 <= 0;
        Res_3_1 <= 0;
        Res_3_2 <= 0;
        Res_3_3 <= 0;
        Res_3_4 <= 0;
        Res_3_5 <= 0;
        Res_3_6 <= 0;
        Res_3_7 <= 0;
        Res_4_0 <= 0;
        Res_4_1 <= 0;
        Res_4_2 <= 0;
        Res_4_3 <= 0;
        Res_4_4 <= 0;
        Res_4_5 <= 0;
        Res_4_6 <= 0;
        Res_4_7 <= 0;
        Res_5_0 <= 0;
        Res_5_1 <= 0;
        Res_5_2 <= 0;
        Res_5_3 <= 0;
        Res_5_4 <= 0;
        Res_5_5 <= 0;
        Res_5_6 <= 0;
        Res_5_7 <= 0;
        Res_6_0 <= 0;
        Res_6_1 <= 0;
        Res_6_2 <= 0;
        Res_6_3 <= 0;
        Res_6_4 <= 0;
        Res_6_5 <= 0;
        Res_6_6 <= 0;
        Res_6_7 <= 0;
        Res_7_0 <= 0;
        Res_7_1 <= 0;
        Res_7_2 <= 0;
        Res_7_3 <= 0;
        Res_7_4 <= 0;
        Res_7_5 <= 0;
        Res_7_6 <= 0;
        Res_7_7 <= 0;
        Res_8_0 <= 0;
        Res_8_1 <= 0;
        Res_8_2 <= 0;
        Res_8_3 <= 0;
        Res_8_4 <= 0;
        Res_8_5 <= 0;
        Res_8_6 <= 0;
        Res_8_7 <= 0;
        Res_9_0 <= 0;
        Res_9_1 <= 0;
        Res_9_2 <= 0;
        Res_9_3 <= 0;
        Res_9_4 <= 0;
        Res_9_5 <= 0;
        Res_9_6 <= 0;
        Res_9_7 <= 0;

    end
    else begin
        Res_0_0<= Res_0_0_n;
        Res_0_1<= Res_0_1_n;
        Res_0_2<= Res_0_2_n;
        Res_0_3<= Res_0_3_n;
        Res_0_4<= Res_0_4_n;
        Res_0_5<= Res_0_5_n;
        Res_0_6<= Res_0_6_n;
        Res_0_7<= Res_0_7_n;
        Res_1_0<= Res_1_0_n;
        Res_1_1<= Res_1_1_n;
        Res_1_2<= Res_1_2_n;
        Res_1_3<= Res_1_3_n;
        Res_1_4<= Res_1_4_n;
        Res_1_5<= Res_1_5_n;
        Res_1_6<= Res_1_6_n;
        Res_1_7<= Res_1_7_n;
        Res_2_0<= Res_2_0_n;
        Res_2_1<= Res_2_1_n;
        Res_2_2<= Res_2_2_n;
        Res_2_3<= Res_2_3_n;
        Res_2_4<= Res_2_4_n;
        Res_2_5<= Res_2_5_n;
        Res_2_6<= Res_2_6_n;
        Res_2_7<= Res_2_7_n;
        Res_3_0<= Res_3_0_n;
        Res_3_1<= Res_3_1_n;
        Res_3_2<= Res_3_2_n;
        Res_3_3<= Res_3_3_n;
        Res_3_4<= Res_3_4_n;
        Res_3_5<= Res_3_5_n;
        Res_3_6<= Res_3_6_n;
        Res_3_7<= Res_3_7_n;
        Res_4_0<= Res_4_0_n;
        Res_4_1<= Res_4_1_n;
        Res_4_2<= Res_4_2_n;
        Res_4_3<= Res_4_3_n;
        Res_4_4<= Res_4_4_n;
        Res_4_5<= Res_4_5_n;
        Res_4_6<= Res_4_6_n;
        Res_4_7<= Res_4_7_n;
        Res_5_0<= Res_5_0_n;
        Res_5_1<= Res_5_1_n;
        Res_5_2<= Res_5_2_n;
        Res_5_3<= Res_5_3_n;
        Res_5_4<= Res_5_4_n;
        Res_5_5<= Res_5_5_n;
        Res_5_6<= Res_5_6_n;
        Res_5_7<= Res_5_7_n;
        Res_6_0<= Res_6_0_n;
        Res_6_1<= Res_6_1_n;
        Res_6_2<= Res_6_2_n;
        Res_6_3<= Res_6_3_n;
        Res_6_4<= Res_6_4_n;
        Res_6_5<= Res_6_5_n;
        Res_6_6<= Res_6_6_n;
        Res_6_7<= Res_6_7_n;
        Res_7_0<= Res_7_0_n;
        Res_7_1<= Res_7_1_n;
        Res_7_2<= Res_7_2_n;
        Res_7_3<= Res_7_3_n;
        Res_7_4<= Res_7_4_n;
        Res_7_5<= Res_7_5_n;
        Res_7_6<= Res_7_6_n;
        Res_7_7<= Res_7_7_n;
        Res_8_0<= Res_8_0_n;
        Res_8_1<= Res_8_1_n;
        Res_8_2<= Res_8_2_n;
        Res_8_3<= Res_8_3_n;
        Res_8_4<= Res_8_4_n;
        Res_8_5<= Res_8_5_n;
        Res_8_6<= Res_8_6_n;
        Res_8_7<= Res_8_7_n;
        Res_9_0<= Res_9_0_n;
        Res_9_1<= Res_9_1_n;
        Res_9_2<= Res_9_2_n;
        Res_9_3<= Res_9_3_n;
        Res_9_4<= Res_9_4_n;
        Res_9_5<= Res_9_5_n;
        Res_9_6<= Res_9_6_n;
        Res_9_7<= Res_9_7_n;

    end
end

// Result assignment
assign Image_Number = V31>V32? W31:W32;
/////////////////////////////////////////////////////////
// Generate blocks
// Registers inside Multipler
generate
genvar a;
for(a=0; a<784/8; a=a+1)begin: Mult_Buf
    reg [9:0]  Feature;
    reg [18:0] Weight;
    reg [9:0]  Feature_n;
    reg [18:0] Weight_n;
    always@(posedge clk, negedge GlobalReset)begin
        if(!GlobalReset)begin
            Weight <=0;
            Feature <=0;
        end
        else begin
            Weight <= Weight_n;
            Feature<=Feature_n;
        end
    end
end
endgenerate

// Registers inside adders
generate
genvar b;
for(b=0; b<49; b=b+1)begin: Add_Buf
    reg[25:0]  A;
    reg[25:0]  B;
    reg[25:0]  A_n;
    reg[25:0]  B_n;
    always@(posedge clk, negedge GlobalReset)begin
        if(!GlobalReset)begin
            A <=0;
            B <=0;
        end
        else begin
            A <= A_n;
            B <= B_n;
        end
    end
end
endgenerate
//////// Multiplier Instantiation///////
genvar i;
// Instantiate 0-195 Mutiplyer
generate
for (i=0; i<784/8; i = i+1) begin: Multiplyer_matrix
    wire[25:0] Result;
    FixedPointMultiplier Inst(.clk(clk),.GlobalReset(~GlobalReset),.WeightPort(Mult_Buf[i].Weight),.PixelPort(Mult_Buf[i].Feature[8:0]),.Output_syn(Result));
end
endgenerate
// Instantiate 6 level Adder Tree, total dealy = 14; Partially TESTED
    wire[25:0] Part_Res;
    wire[25:0] Final_Res;
    // Base
    // L1
    
    genvar k;
    generate
    for(k = 0; k<49; k=k+1) begin:Adder_Base
        wire[25:0] Res;
        FixedPointAdder Adder( .clk(clk),.GlobalReset(~GlobalReset),.Port1(Add_Buf[k].A),.Port2(Add_Buf[k].B),.Output_syn(Res));
    end
    endgenerate

    // L2
    genvar l;
    generate
    for(l=0; l<25; l=l+1) begin:Adder_L2
        wire[25:0] Res;
        if(l<24)
            FixedPointAdder Adder( .clk(clk),.GlobalReset(~GlobalReset),.Port1(Adder_Base[l*2].Res),.Port2(Adder_Base[l*2+1].Res),.Output_syn(Res));
        else
            FixedPointAdder Adder( .clk(clk),.GlobalReset(~GlobalReset),.Port1(Adder_Base[l*2].Res),.Port2(26'b0),.Output_syn(Res));
    end
    endgenerate

    // L3
    genvar m;
    generate
    for(m=0; m<13; m=m+1) begin:Adder_L3
        wire[25:0] Res;
        if(m<12)
            FixedPointAdder Adder( .clk(clk),.GlobalReset(~GlobalReset),.Port1(Adder_L2[m*2].Res),.Port2(Adder_L2[m*2+1].Res),.Output_syn(Res));
        else
            FixedPointAdder Adder( .clk(clk),.GlobalReset(~GlobalReset),.Port1(Adder_L2[m*2].Res),.Port2(26'b0),.Output_syn(Res));
    end
    endgenerate

    // L4
    genvar n;
    generate
    for(n=0; n<7; n=n+1) begin:Adder_L4
        wire[25:0] Res;
        if(n < 6)
            FixedPointAdder Adder( .clk(clk),.GlobalReset(~GlobalReset),.Port1(Adder_L3[n*2].Res),.Port2(Adder_L3[n*2+1].Res),.Output_syn(Res));
        else 
            FixedPointAdder Adder( .clk(clk),.GlobalReset(~GlobalReset),.Port1(Adder_L3[n*2].Res),.Port2(26'b0),.Output_syn(Res));
    end
    endgenerate

    // L5
    genvar o;
    generate
    for(o=0; o<4; o=o+1) begin:Adder_L5
        wire[25:0] Res;
        if(o < 3)
            FixedPointAdder Adder( .clk(clk),.GlobalReset(~GlobalReset),.Port1(Adder_L4[o*2].Res),.Port2(Adder_L4[o*2+1].Res),.Output_syn(Res));
        else
            FixedPointAdder Adder( .clk(clk),.GlobalReset(~GlobalReset),.Port1(Adder_L4[o*2].Res),.Port2(26'b0),.Output_syn(Res));
    end
    endgenerate

    // L6
    genvar p;
    generate
    for(p=0; p<2;p=p+1) begin:Adder_L6
        wire[25:0] Res;
            FixedPointAdder Adder( .clk(clk),.GlobalReset(~GlobalReset),.Port1(Adder_L5[p*2].Res),.Port2(Adder_L5[p*2+1].Res),.Output_syn(Res));
    end
    endgenerate

    // L7
    FixedPointAdder FinalAdder( .clk(clk),.GlobalReset(~GlobalReset),.Port1(Adder_L6[0].Res),.Port2(Adder_L6[1].Res),.Output_syn(Part_Res));

//////// Instantiate three final adder//////    6 cycle delay
    reg [25:0]A1,A2,A3,A4,A5,A6,A7,A8;
    wire [25:0]B1,B2,B3,B4;
    wire [25:0]C1,C2;

    FixedPointAdder Adder_A1( .clk(clk),.GlobalReset(~GlobalReset),.Port1(A1),.Port2(A2),.Output_syn(B1));
    FixedPointAdder Adder_A3( .clk(clk),.GlobalReset(~GlobalReset),.Port1(A3),.Port2(A4),.Output_syn(B2));
    FixedPointAdder Adder_A5( .clk(clk),.GlobalReset(~GlobalReset),.Port1(A5),.Port2(A6),.Output_syn(B3));
    FixedPointAdder Adder_A6( .clk(clk),.GlobalReset(~GlobalReset),.Port1(A7),.Port2(A8),.Output_syn(B4));

    FixedPointAdder Adder_B1( .clk(clk),.GlobalReset(~GlobalReset),.Port1(B1),.Port2(B2),.Output_syn(C1));
    FixedPointAdder Adder_B2( .clk(clk),.GlobalReset(~GlobalReset),.Port1(B3),.Port2(B4),.Output_syn(C2));

    FixedPointAdder Top( .clk(clk),.GlobalReset(~GlobalReset),.Port1(C1),.Port2(C2),.Output_syn(Final_Res));

//////// State Transition Logic///////////
always@(*)begin
    Load = 0;
    nxt_state = 0;
    Add_Buf[0].A_n = 0;
        Add_Buf[0].B_n = 0;
        Add_Buf[1].A_n = 0;
        Add_Buf[1].B_n = 0;
        Add_Buf[2].A_n = 0;
        Add_Buf[2].B_n = 0;
        Add_Buf[3].A_n = 0;
        Add_Buf[3].B_n = 0;
        Add_Buf[4].A_n = 0;
        Add_Buf[4].B_n = 0;
        Add_Buf[5].A_n = 0;
        Add_Buf[5].B_n = 0;
        Add_Buf[6].A_n = 0;
        Add_Buf[6].B_n = 0;
        Add_Buf[7].A_n = 0;
        Add_Buf[7].B_n = 0;
        Add_Buf[8].A_n = 0;
        Add_Buf[8].B_n = 0;
        Add_Buf[9].A_n = 0;
        Add_Buf[9].B_n = 0;
        Add_Buf[10].A_n = 0;
        Add_Buf[10].B_n = 0;
        Add_Buf[11].A_n = 0;
        Add_Buf[11].B_n = 0;
        Add_Buf[12].A_n = 0;
        Add_Buf[12].B_n = 0;
        Add_Buf[13].A_n = 0;
        Add_Buf[13].B_n = 0;
        Add_Buf[14].A_n = 0;
        Add_Buf[14].B_n = 0;
        Add_Buf[15].A_n = 0;
        Add_Buf[15].B_n = 0;
        Add_Buf[16].A_n = 0;
        Add_Buf[16].B_n = 0;
        Add_Buf[17].A_n = 0;
        Add_Buf[17].B_n = 0;
        Add_Buf[18].A_n = 0;
        Add_Buf[18].B_n = 0;
        Add_Buf[19].A_n = 0;
        Add_Buf[19].B_n = 0;
        Add_Buf[20].A_n = 0;
        Add_Buf[20].B_n = 0;
        Add_Buf[21].A_n = 0;
        Add_Buf[21].B_n = 0;
        Add_Buf[22].A_n = 0;
        Add_Buf[22].B_n = 0;
        Add_Buf[23].A_n = 0;
        Add_Buf[23].B_n = 0;
        Add_Buf[24].A_n = 0;
        Add_Buf[24].B_n = 0;
        Add_Buf[25].A_n = 0;
        Add_Buf[25].B_n = 0;
        Add_Buf[26].A_n = 0;
        Add_Buf[26].B_n = 0;
        Add_Buf[27].A_n = 0;
        Add_Buf[27].B_n = 0;
        Add_Buf[28].A_n = 0;
        Add_Buf[28].B_n = 0;
        Add_Buf[29].A_n = 0;
        Add_Buf[29].B_n = 0;
        Add_Buf[30].A_n = 0;
        Add_Buf[30].B_n = 0;
        Add_Buf[31].A_n = 0;
        Add_Buf[31].B_n = 0;
        Add_Buf[32].A_n = 0;
        Add_Buf[32].B_n = 0;
        Add_Buf[33].A_n = 0;
        Add_Buf[33].B_n = 0;
        Add_Buf[34].A_n = 0;
        Add_Buf[34].B_n = 0;
        Add_Buf[35].A_n = 0;
        Add_Buf[35].B_n = 0;
        Add_Buf[36].A_n = 0;
        Add_Buf[36].B_n = 0;
        Add_Buf[37].A_n = 0;
        Add_Buf[37].B_n = 0;
        Add_Buf[38].A_n = 0;
        Add_Buf[38].B_n = 0;
        Add_Buf[39].A_n = 0;
        Add_Buf[39].B_n = 0;
        Add_Buf[40].A_n = 0;
        Add_Buf[40].B_n = 0;
        Add_Buf[41].A_n = 0;
        Add_Buf[41].B_n = 0;
        Add_Buf[42].A_n = 0;
        Add_Buf[42].B_n = 0;
        Add_Buf[43].A_n = 0;
        Add_Buf[43].B_n = 0;
        Add_Buf[44].A_n = 0;
        Add_Buf[44].B_n = 0;
        Add_Buf[45].A_n = 0;
        Add_Buf[45].B_n = 0;
        Add_Buf[46].A_n = 0;
        Add_Buf[46].B_n = 0;
        Add_Buf[47].A_n = 0;
        Add_Buf[47].B_n = 0;
        Add_Buf[48].A_n = 0;
        Add_Buf[48].B_n = 0;

    Mult_Buf[0].Weight_n = 0;
        Mult_Buf[0].Feature_n = 0;
        Mult_Buf[1].Weight_n = 0;
        Mult_Buf[1].Feature_n = 0;
        Mult_Buf[2].Weight_n = 0;
        Mult_Buf[2].Feature_n = 0;
        Mult_Buf[3].Weight_n = 0;
        Mult_Buf[3].Feature_n = 0;
        Mult_Buf[4].Weight_n = 0;
        Mult_Buf[4].Feature_n = 0;
        Mult_Buf[5].Weight_n = 0;
        Mult_Buf[5].Feature_n = 0;
        Mult_Buf[6].Weight_n = 0;
        Mult_Buf[6].Feature_n = 0;
        Mult_Buf[7].Weight_n = 0;
        Mult_Buf[7].Feature_n = 0;
        Mult_Buf[8].Weight_n = 0;
        Mult_Buf[8].Feature_n = 0;
        Mult_Buf[9].Weight_n = 0;
        Mult_Buf[9].Feature_n = 0;
        Mult_Buf[10].Weight_n = 0;
        Mult_Buf[10].Feature_n = 0;
        Mult_Buf[11].Weight_n = 0;
        Mult_Buf[11].Feature_n = 0;
        Mult_Buf[12].Weight_n = 0;
        Mult_Buf[12].Feature_n = 0;
        Mult_Buf[13].Weight_n = 0;
        Mult_Buf[13].Feature_n = 0;
        Mult_Buf[14].Weight_n = 0;
        Mult_Buf[14].Feature_n = 0;
        Mult_Buf[15].Weight_n = 0;
        Mult_Buf[15].Feature_n = 0;
        Mult_Buf[16].Weight_n = 0;
        Mult_Buf[16].Feature_n = 0;
        Mult_Buf[17].Weight_n = 0;
        Mult_Buf[17].Feature_n = 0;
        Mult_Buf[18].Weight_n = 0;
        Mult_Buf[18].Feature_n = 0;
        Mult_Buf[19].Weight_n = 0;
        Mult_Buf[19].Feature_n = 0;
        Mult_Buf[20].Weight_n = 0;
        Mult_Buf[20].Feature_n = 0;
        Mult_Buf[21].Weight_n = 0;
        Mult_Buf[21].Feature_n = 0;
        Mult_Buf[22].Weight_n = 0;
        Mult_Buf[22].Feature_n = 0;
        Mult_Buf[23].Weight_n = 0;
        Mult_Buf[23].Feature_n = 0;
        Mult_Buf[24].Weight_n = 0;
        Mult_Buf[24].Feature_n = 0;
        Mult_Buf[25].Weight_n = 0;
        Mult_Buf[25].Feature_n = 0;
        Mult_Buf[26].Weight_n = 0;
        Mult_Buf[26].Feature_n = 0;
        Mult_Buf[27].Weight_n = 0;
        Mult_Buf[27].Feature_n = 0;
        Mult_Buf[28].Weight_n = 0;
        Mult_Buf[28].Feature_n = 0;
        Mult_Buf[29].Weight_n = 0;
        Mult_Buf[29].Feature_n = 0;
        Mult_Buf[30].Weight_n = 0;
        Mult_Buf[30].Feature_n = 0;
        Mult_Buf[31].Weight_n = 0;
        Mult_Buf[31].Feature_n = 0;
        Mult_Buf[32].Weight_n = 0;
        Mult_Buf[32].Feature_n = 0;
        Mult_Buf[33].Weight_n = 0;
        Mult_Buf[33].Feature_n = 0;
        Mult_Buf[34].Weight_n = 0;
        Mult_Buf[34].Feature_n = 0;
        Mult_Buf[35].Weight_n = 0;
        Mult_Buf[35].Feature_n = 0;
        Mult_Buf[36].Weight_n = 0;
        Mult_Buf[36].Feature_n = 0;
        Mult_Buf[37].Weight_n = 0;
        Mult_Buf[37].Feature_n = 0;
        Mult_Buf[38].Weight_n = 0;
        Mult_Buf[38].Feature_n = 0;
        Mult_Buf[39].Weight_n = 0;
        Mult_Buf[39].Feature_n = 0;
        Mult_Buf[40].Weight_n = 0;
        Mult_Buf[40].Feature_n = 0;
        Mult_Buf[41].Weight_n = 0;
        Mult_Buf[41].Feature_n = 0;
        Mult_Buf[42].Weight_n = 0;
        Mult_Buf[42].Feature_n = 0;
        Mult_Buf[43].Weight_n = 0;
        Mult_Buf[43].Feature_n = 0;
        Mult_Buf[44].Weight_n = 0;
        Mult_Buf[44].Feature_n = 0;
        Mult_Buf[45].Weight_n = 0;
        Mult_Buf[45].Feature_n = 0;
        Mult_Buf[46].Weight_n = 0;
        Mult_Buf[46].Feature_n = 0;
        Mult_Buf[47].Weight_n = 0;
        Mult_Buf[47].Feature_n = 0;
        Mult_Buf[48].Weight_n = 0;
        Mult_Buf[48].Feature_n = 0;
        Mult_Buf[49].Weight_n = 0;
        Mult_Buf[49].Feature_n = 0;
        Mult_Buf[50].Weight_n = 0;
        Mult_Buf[50].Feature_n = 0;
        Mult_Buf[51].Weight_n = 0;
        Mult_Buf[51].Feature_n = 0;
        Mult_Buf[52].Weight_n = 0;
        Mult_Buf[52].Feature_n = 0;
        Mult_Buf[53].Weight_n = 0;
        Mult_Buf[53].Feature_n = 0;
        Mult_Buf[54].Weight_n = 0;
        Mult_Buf[54].Feature_n = 0;
        Mult_Buf[55].Weight_n = 0;
        Mult_Buf[55].Feature_n = 0;
        Mult_Buf[56].Weight_n = 0;
        Mult_Buf[56].Feature_n = 0;
        Mult_Buf[57].Weight_n = 0;
        Mult_Buf[57].Feature_n = 0;
        Mult_Buf[58].Weight_n = 0;
        Mult_Buf[58].Feature_n = 0;
        Mult_Buf[59].Weight_n = 0;
        Mult_Buf[59].Feature_n = 0;
        Mult_Buf[60].Weight_n = 0;
        Mult_Buf[60].Feature_n = 0;
        Mult_Buf[61].Weight_n = 0;
        Mult_Buf[61].Feature_n = 0;
        Mult_Buf[62].Weight_n = 0;
        Mult_Buf[62].Feature_n = 0;
        Mult_Buf[63].Weight_n = 0;
        Mult_Buf[63].Feature_n = 0;
        Mult_Buf[64].Weight_n = 0;
        Mult_Buf[64].Feature_n = 0;
        Mult_Buf[65].Weight_n = 0;
        Mult_Buf[65].Feature_n = 0;
        Mult_Buf[66].Weight_n = 0;
        Mult_Buf[66].Feature_n = 0;
        Mult_Buf[67].Weight_n = 0;
        Mult_Buf[67].Feature_n = 0;
        Mult_Buf[68].Weight_n = 0;
        Mult_Buf[68].Feature_n = 0;
        Mult_Buf[69].Weight_n = 0;
        Mult_Buf[69].Feature_n = 0;
        Mult_Buf[70].Weight_n = 0;
        Mult_Buf[70].Feature_n = 0;
        Mult_Buf[71].Weight_n = 0;
        Mult_Buf[71].Feature_n = 0;
        Mult_Buf[72].Weight_n = 0;
        Mult_Buf[72].Feature_n = 0;
        Mult_Buf[73].Weight_n = 0;
        Mult_Buf[73].Feature_n = 0;
        Mult_Buf[74].Weight_n = 0;
        Mult_Buf[74].Feature_n = 0;
        Mult_Buf[75].Weight_n = 0;
        Mult_Buf[75].Feature_n = 0;
        Mult_Buf[76].Weight_n = 0;
        Mult_Buf[76].Feature_n = 0;
        Mult_Buf[77].Weight_n = 0;
        Mult_Buf[77].Feature_n = 0;
        Mult_Buf[78].Weight_n = 0;
        Mult_Buf[78].Feature_n = 0;
        Mult_Buf[79].Weight_n = 0;
        Mult_Buf[79].Feature_n = 0;
        Mult_Buf[80].Weight_n = 0;
        Mult_Buf[80].Feature_n = 0;
        Mult_Buf[81].Weight_n = 0;
        Mult_Buf[81].Feature_n = 0;
        Mult_Buf[82].Weight_n = 0;
        Mult_Buf[82].Feature_n = 0;
        Mult_Buf[83].Weight_n = 0;
        Mult_Buf[83].Feature_n = 0;
        Mult_Buf[84].Weight_n = 0;
        Mult_Buf[84].Feature_n = 0;
        Mult_Buf[85].Weight_n = 0;
        Mult_Buf[85].Feature_n = 0;
        Mult_Buf[86].Weight_n = 0;
        Mult_Buf[86].Feature_n = 0;
        Mult_Buf[87].Weight_n = 0;
        Mult_Buf[87].Feature_n = 0;
        Mult_Buf[88].Weight_n = 0;
        Mult_Buf[88].Feature_n = 0;
        Mult_Buf[89].Weight_n = 0;
        Mult_Buf[89].Feature_n = 0;
        Mult_Buf[90].Weight_n = 0;
        Mult_Buf[90].Feature_n = 0;
        Mult_Buf[91].Weight_n = 0;
        Mult_Buf[91].Feature_n = 0;
        Mult_Buf[92].Weight_n = 0;
        Mult_Buf[92].Feature_n = 0;
        Mult_Buf[93].Weight_n = 0;
        Mult_Buf[93].Feature_n = 0;
        Mult_Buf[94].Weight_n = 0;
        Mult_Buf[94].Feature_n = 0;
        Mult_Buf[95].Weight_n = 0;
        Mult_Buf[95].Feature_n = 0;
        Mult_Buf[96].Weight_n = 0;
        Mult_Buf[96].Feature_n = 0;
        Mult_Buf[97].Weight_n = 0;
        Mult_Buf[97].Feature_n = 0;


    Res_0_0_n = Res_0_0;
        Res_0_1_n = Res_0_1;
        Res_0_2_n = Res_0_2;
        Res_0_3_n = Res_0_3;
        Res_0_4_n = Res_0_4;
        Res_0_5_n = Res_0_5;
        Res_0_6_n = Res_0_6;
        Res_0_7_n = Res_0_7;
        Res_1_0_n = Res_1_0;
        Res_1_1_n = Res_1_1;
        Res_1_2_n = Res_1_2;
        Res_1_3_n = Res_1_3;
        Res_1_4_n = Res_1_4;
        Res_1_5_n = Res_1_5;
        Res_1_6_n = Res_1_6;
        Res_1_7_n = Res_1_7;
        Res_2_0_n = Res_2_0;
        Res_2_1_n = Res_2_1;
        Res_2_2_n = Res_2_2;
        Res_2_3_n = Res_2_3;
        Res_2_4_n = Res_2_4;
        Res_2_5_n = Res_2_5;
        Res_2_6_n = Res_2_6;
        Res_2_7_n = Res_2_7;
        Res_3_0_n = Res_3_0;
        Res_3_1_n = Res_3_1;
        Res_3_2_n = Res_3_2;
        Res_3_3_n = Res_3_3;
        Res_3_4_n = Res_3_4;
        Res_3_5_n = Res_3_5;
        Res_3_6_n = Res_3_6;
        Res_3_7_n = Res_3_7;
        Res_4_0_n = Res_4_0;
        Res_4_1_n = Res_4_1;
        Res_4_2_n = Res_4_2;
        Res_4_3_n = Res_4_3;
        Res_4_4_n = Res_4_4;
        Res_4_5_n = Res_4_5;
        Res_4_6_n = Res_4_6;
        Res_4_7_n = Res_4_7;
        Res_5_0_n = Res_5_0;
        Res_5_1_n = Res_5_1;
        Res_5_2_n = Res_5_2;
        Res_5_3_n = Res_5_3;
        Res_5_4_n = Res_5_4;
        Res_5_5_n = Res_5_5;
        Res_5_6_n = Res_5_6;
        Res_5_7_n = Res_5_7;
        Res_6_0_n = Res_6_0;
        Res_6_1_n = Res_6_1;
        Res_6_2_n = Res_6_2;
        Res_6_3_n = Res_6_3;
        Res_6_4_n = Res_6_4;
        Res_6_5_n = Res_6_5;
        Res_6_6_n = Res_6_6;
        Res_6_7_n = Res_6_7;
        Res_7_0_n = Res_7_0;
        Res_7_1_n = Res_7_1;
        Res_7_2_n = Res_7_2;
        Res_7_3_n = Res_7_3;
        Res_7_4_n = Res_7_4;
        Res_7_5_n = Res_7_5;
        Res_7_6_n = Res_7_6;
        Res_7_7_n = Res_7_7;
        Res_8_0_n = Res_8_0;
        Res_8_1_n = Res_8_1;
        Res_8_2_n = Res_8_2;
        Res_8_3_n = Res_8_3;
        Res_8_4_n = Res_8_4;
        Res_8_5_n = Res_8_5;
        Res_8_6_n = Res_8_6;
        Res_8_7_n = Res_8_7;
        Res_9_0_n = Res_9_0;
        Res_9_1_n = Res_9_1;
        Res_9_2_n = Res_9_2;
        Res_9_3_n = Res_9_3;
        Res_9_4_n = Res_9_4;
        Res_9_5_n = Res_9_5;
        Res_9_6_n = Res_9_6;
        Res_9_7_n = Res_9_7;


    Res0_n = Res0;
        Res1_n = Res1;
        Res2_n = Res2;
        Res3_n = Res3;
        Res4_n = Res4;
        Res5_n = Res5;
        Res6_n = Res6;
        Res7_n = Res7;
        Res8_n = Res8;
        Res9_n = Res9;
    Output_Valid = 0;
      //Initialize value
    A1=0;
        A2=0;
        A3=0;
        A4=0;
        A5=0;
        A6=0;
        A7=0;
        A8=0;
    W11_n = 0;
        W12_n = 0;
        W13_n = 0;
        W14_n = 0;
        W15_n = 0;
        V11_n = 0;
        V12_n = 0;
        V13_n = 0;
        V14_n = 0;
        V15_n = 0;
        W21_n = 0;
        W22_n = 0;
        V21_n = 0;
        V22_n = 0;
        W31_n = 0;
        W32_n = 0;
        V31_n = 0;
        V32_n = 0;
 
    //Ending Initialize value
    case(state)
    // IDLE State
    0:begin
        nxt_state = Input_Valid?1:0;
        end
    // Buffer All Input
    1:begin
        Load = 1;
        nxt_state = 2;
        end
    
   
   

///////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////

    2:begin
     nxt_state = 3;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_0;
         Mult_Buf[0].Weight_n = Wgt_0_0;
         Mult_Buf[1].Feature_n = FeatureBuf_1;
         Mult_Buf[1].Weight_n = Wgt_0_1;
         Mult_Buf[2].Feature_n = FeatureBuf_2;
         Mult_Buf[2].Weight_n = Wgt_0_2;
         Mult_Buf[3].Feature_n = FeatureBuf_3;
         Mult_Buf[3].Weight_n = Wgt_0_3;
         Mult_Buf[4].Feature_n = FeatureBuf_4;
         Mult_Buf[4].Weight_n = Wgt_0_4;
         Mult_Buf[5].Feature_n = FeatureBuf_5;
         Mult_Buf[5].Weight_n = Wgt_0_5;
         Mult_Buf[6].Feature_n = FeatureBuf_6;
         Mult_Buf[6].Weight_n = Wgt_0_6;
         Mult_Buf[7].Feature_n = FeatureBuf_7;
         Mult_Buf[7].Weight_n = Wgt_0_7;
         Mult_Buf[8].Feature_n = FeatureBuf_8;
         Mult_Buf[8].Weight_n = Wgt_0_8;
         Mult_Buf[9].Feature_n = FeatureBuf_9;
         Mult_Buf[9].Weight_n = Wgt_0_9;
         Mult_Buf[10].Feature_n = FeatureBuf_10;
         Mult_Buf[10].Weight_n = Wgt_0_10;
         Mult_Buf[11].Feature_n = FeatureBuf_11;
         Mult_Buf[11].Weight_n = Wgt_0_11;
         Mult_Buf[12].Feature_n = FeatureBuf_12;
         Mult_Buf[12].Weight_n = Wgt_0_12;
         Mult_Buf[13].Feature_n = FeatureBuf_13;
         Mult_Buf[13].Weight_n = Wgt_0_13;
         Mult_Buf[14].Feature_n = FeatureBuf_14;
         Mult_Buf[14].Weight_n = Wgt_0_14;
         Mult_Buf[15].Feature_n = FeatureBuf_15;
         Mult_Buf[15].Weight_n = Wgt_0_15;
         Mult_Buf[16].Feature_n = FeatureBuf_16;
         Mult_Buf[16].Weight_n = Wgt_0_16;
         Mult_Buf[17].Feature_n = FeatureBuf_17;
         Mult_Buf[17].Weight_n = Wgt_0_17;
         Mult_Buf[18].Feature_n = FeatureBuf_18;
         Mult_Buf[18].Weight_n = Wgt_0_18;
         Mult_Buf[19].Feature_n = FeatureBuf_19;
         Mult_Buf[19].Weight_n = Wgt_0_19;
         Mult_Buf[20].Feature_n = FeatureBuf_20;
         Mult_Buf[20].Weight_n = Wgt_0_20;
         Mult_Buf[21].Feature_n = FeatureBuf_21;
         Mult_Buf[21].Weight_n = Wgt_0_21;
         Mult_Buf[22].Feature_n = FeatureBuf_22;
         Mult_Buf[22].Weight_n = Wgt_0_22;
         Mult_Buf[23].Feature_n = FeatureBuf_23;
         Mult_Buf[23].Weight_n = Wgt_0_23;
         Mult_Buf[24].Feature_n = FeatureBuf_24;
         Mult_Buf[24].Weight_n = Wgt_0_24;
         Mult_Buf[25].Feature_n = FeatureBuf_25;
         Mult_Buf[25].Weight_n = Wgt_0_25;
         Mult_Buf[26].Feature_n = FeatureBuf_26;
         Mult_Buf[26].Weight_n = Wgt_0_26;
         Mult_Buf[27].Feature_n = FeatureBuf_27;
         Mult_Buf[27].Weight_n = Wgt_0_27;
         Mult_Buf[28].Feature_n = FeatureBuf_28;
         Mult_Buf[28].Weight_n = Wgt_0_28;
         Mult_Buf[29].Feature_n = FeatureBuf_29;
         Mult_Buf[29].Weight_n = Wgt_0_29;
         Mult_Buf[30].Feature_n = FeatureBuf_30;
         Mult_Buf[30].Weight_n = Wgt_0_30;
         Mult_Buf[31].Feature_n = FeatureBuf_31;
         Mult_Buf[31].Weight_n = Wgt_0_31;
         Mult_Buf[32].Feature_n = FeatureBuf_32;
         Mult_Buf[32].Weight_n = Wgt_0_32;
         Mult_Buf[33].Feature_n = FeatureBuf_33;
         Mult_Buf[33].Weight_n = Wgt_0_33;
         Mult_Buf[34].Feature_n = FeatureBuf_34;
         Mult_Buf[34].Weight_n = Wgt_0_34;
         Mult_Buf[35].Feature_n = FeatureBuf_35;
         Mult_Buf[35].Weight_n = Wgt_0_35;
         Mult_Buf[36].Feature_n = FeatureBuf_36;
         Mult_Buf[36].Weight_n = Wgt_0_36;
         Mult_Buf[37].Feature_n = FeatureBuf_37;
         Mult_Buf[37].Weight_n = Wgt_0_37;
         Mult_Buf[38].Feature_n = FeatureBuf_38;
         Mult_Buf[38].Weight_n = Wgt_0_38;
         Mult_Buf[39].Feature_n = FeatureBuf_39;
         Mult_Buf[39].Weight_n = Wgt_0_39;
         Mult_Buf[40].Feature_n = FeatureBuf_40;
         Mult_Buf[40].Weight_n = Wgt_0_40;
         Mult_Buf[41].Feature_n = FeatureBuf_41;
         Mult_Buf[41].Weight_n = Wgt_0_41;
         Mult_Buf[42].Feature_n = FeatureBuf_42;
         Mult_Buf[42].Weight_n = Wgt_0_42;
         Mult_Buf[43].Feature_n = FeatureBuf_43;
         Mult_Buf[43].Weight_n = Wgt_0_43;
         Mult_Buf[44].Feature_n = FeatureBuf_44;
         Mult_Buf[44].Weight_n = Wgt_0_44;
         Mult_Buf[45].Feature_n = FeatureBuf_45;
         Mult_Buf[45].Weight_n = Wgt_0_45;
         Mult_Buf[46].Feature_n = FeatureBuf_46;
         Mult_Buf[46].Weight_n = Wgt_0_46;
         Mult_Buf[47].Feature_n = FeatureBuf_47;
         Mult_Buf[47].Weight_n = Wgt_0_47;
         Mult_Buf[48].Feature_n = FeatureBuf_48;
         Mult_Buf[48].Weight_n = Wgt_0_48;
         Mult_Buf[49].Feature_n = FeatureBuf_49;
         Mult_Buf[49].Weight_n = Wgt_0_49;
         Mult_Buf[50].Feature_n = FeatureBuf_50;
         Mult_Buf[50].Weight_n = Wgt_0_50;
         Mult_Buf[51].Feature_n = FeatureBuf_51;
         Mult_Buf[51].Weight_n = Wgt_0_51;
         Mult_Buf[52].Feature_n = FeatureBuf_52;
         Mult_Buf[52].Weight_n = Wgt_0_52;
         Mult_Buf[53].Feature_n = FeatureBuf_53;
         Mult_Buf[53].Weight_n = Wgt_0_53;
         Mult_Buf[54].Feature_n = FeatureBuf_54;
         Mult_Buf[54].Weight_n = Wgt_0_54;
         Mult_Buf[55].Feature_n = FeatureBuf_55;
         Mult_Buf[55].Weight_n = Wgt_0_55;
         Mult_Buf[56].Feature_n = FeatureBuf_56;
         Mult_Buf[56].Weight_n = Wgt_0_56;
         Mult_Buf[57].Feature_n = FeatureBuf_57;
         Mult_Buf[57].Weight_n = Wgt_0_57;
         Mult_Buf[58].Feature_n = FeatureBuf_58;
         Mult_Buf[58].Weight_n = Wgt_0_58;
         Mult_Buf[59].Feature_n = FeatureBuf_59;
         Mult_Buf[59].Weight_n = Wgt_0_59;
         Mult_Buf[60].Feature_n = FeatureBuf_60;
         Mult_Buf[60].Weight_n = Wgt_0_60;
         Mult_Buf[61].Feature_n = FeatureBuf_61;
         Mult_Buf[61].Weight_n = Wgt_0_61;
         Mult_Buf[62].Feature_n = FeatureBuf_62;
         Mult_Buf[62].Weight_n = Wgt_0_62;
         Mult_Buf[63].Feature_n = FeatureBuf_63;
         Mult_Buf[63].Weight_n = Wgt_0_63;
         Mult_Buf[64].Feature_n = FeatureBuf_64;
         Mult_Buf[64].Weight_n = Wgt_0_64;
         Mult_Buf[65].Feature_n = FeatureBuf_65;
         Mult_Buf[65].Weight_n = Wgt_0_65;
         Mult_Buf[66].Feature_n = FeatureBuf_66;
         Mult_Buf[66].Weight_n = Wgt_0_66;
         Mult_Buf[67].Feature_n = FeatureBuf_67;
         Mult_Buf[67].Weight_n = Wgt_0_67;
         Mult_Buf[68].Feature_n = FeatureBuf_68;
         Mult_Buf[68].Weight_n = Wgt_0_68;
         Mult_Buf[69].Feature_n = FeatureBuf_69;
         Mult_Buf[69].Weight_n = Wgt_0_69;
         Mult_Buf[70].Feature_n = FeatureBuf_70;
         Mult_Buf[70].Weight_n = Wgt_0_70;
         Mult_Buf[71].Feature_n = FeatureBuf_71;
         Mult_Buf[71].Weight_n = Wgt_0_71;
         Mult_Buf[72].Feature_n = FeatureBuf_72;
         Mult_Buf[72].Weight_n = Wgt_0_72;
         Mult_Buf[73].Feature_n = FeatureBuf_73;
         Mult_Buf[73].Weight_n = Wgt_0_73;
         Mult_Buf[74].Feature_n = FeatureBuf_74;
         Mult_Buf[74].Weight_n = Wgt_0_74;
         Mult_Buf[75].Feature_n = FeatureBuf_75;
         Mult_Buf[75].Weight_n = Wgt_0_75;
         Mult_Buf[76].Feature_n = FeatureBuf_76;
         Mult_Buf[76].Weight_n = Wgt_0_76;
         Mult_Buf[77].Feature_n = FeatureBuf_77;
         Mult_Buf[77].Weight_n = Wgt_0_77;
         Mult_Buf[78].Feature_n = FeatureBuf_78;
         Mult_Buf[78].Weight_n = Wgt_0_78;
         Mult_Buf[79].Feature_n = FeatureBuf_79;
         Mult_Buf[79].Weight_n = Wgt_0_79;
         Mult_Buf[80].Feature_n = FeatureBuf_80;
         Mult_Buf[80].Weight_n = Wgt_0_80;
         Mult_Buf[81].Feature_n = FeatureBuf_81;
         Mult_Buf[81].Weight_n = Wgt_0_81;
         Mult_Buf[82].Feature_n = FeatureBuf_82;
         Mult_Buf[82].Weight_n = Wgt_0_82;
         Mult_Buf[83].Feature_n = FeatureBuf_83;
         Mult_Buf[83].Weight_n = Wgt_0_83;
         Mult_Buf[84].Feature_n = FeatureBuf_84;
         Mult_Buf[84].Weight_n = Wgt_0_84;
         Mult_Buf[85].Feature_n = FeatureBuf_85;
         Mult_Buf[85].Weight_n = Wgt_0_85;
         Mult_Buf[86].Feature_n = FeatureBuf_86;
         Mult_Buf[86].Weight_n = Wgt_0_86;
         Mult_Buf[87].Feature_n = FeatureBuf_87;
         Mult_Buf[87].Weight_n = Wgt_0_87;
         Mult_Buf[88].Feature_n = FeatureBuf_88;
         Mult_Buf[88].Weight_n = Wgt_0_88;
         Mult_Buf[89].Feature_n = FeatureBuf_89;
         Mult_Buf[89].Weight_n = Wgt_0_89;
         Mult_Buf[90].Feature_n = FeatureBuf_90;
         Mult_Buf[90].Weight_n = Wgt_0_90;
         Mult_Buf[91].Feature_n = FeatureBuf_91;
         Mult_Buf[91].Weight_n = Wgt_0_91;
         Mult_Buf[92].Feature_n = FeatureBuf_92;
         Mult_Buf[92].Weight_n = Wgt_0_92;
         Mult_Buf[93].Feature_n = FeatureBuf_93;
         Mult_Buf[93].Weight_n = Wgt_0_93;
         Mult_Buf[94].Feature_n = FeatureBuf_94;
         Mult_Buf[94].Weight_n = Wgt_0_94;
         Mult_Buf[95].Feature_n = FeatureBuf_95;
         Mult_Buf[95].Weight_n = Wgt_0_95;
         Mult_Buf[96].Feature_n = FeatureBuf_96;
         Mult_Buf[96].Weight_n = Wgt_0_96;
         Mult_Buf[97].Feature_n = FeatureBuf_97;
         Mult_Buf[97].Weight_n = Wgt_0_97;
     end
    3:begin
     nxt_state = 4;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_98;
         Mult_Buf[0].Weight_n = Wgt_0_98;
         Mult_Buf[1].Feature_n = FeatureBuf_99;
         Mult_Buf[1].Weight_n = Wgt_0_99;
         Mult_Buf[2].Feature_n = FeatureBuf_100;
         Mult_Buf[2].Weight_n = Wgt_0_100;
         Mult_Buf[3].Feature_n = FeatureBuf_101;
         Mult_Buf[3].Weight_n = Wgt_0_101;
         Mult_Buf[4].Feature_n = FeatureBuf_102;
         Mult_Buf[4].Weight_n = Wgt_0_102;
         Mult_Buf[5].Feature_n = FeatureBuf_103;
         Mult_Buf[5].Weight_n = Wgt_0_103;
         Mult_Buf[6].Feature_n = FeatureBuf_104;
         Mult_Buf[6].Weight_n = Wgt_0_104;
         Mult_Buf[7].Feature_n = FeatureBuf_105;
         Mult_Buf[7].Weight_n = Wgt_0_105;
         Mult_Buf[8].Feature_n = FeatureBuf_106;
         Mult_Buf[8].Weight_n = Wgt_0_106;
         Mult_Buf[9].Feature_n = FeatureBuf_107;
         Mult_Buf[9].Weight_n = Wgt_0_107;
         Mult_Buf[10].Feature_n = FeatureBuf_108;
         Mult_Buf[10].Weight_n = Wgt_0_108;
         Mult_Buf[11].Feature_n = FeatureBuf_109;
         Mult_Buf[11].Weight_n = Wgt_0_109;
         Mult_Buf[12].Feature_n = FeatureBuf_110;
         Mult_Buf[12].Weight_n = Wgt_0_110;
         Mult_Buf[13].Feature_n = FeatureBuf_111;
         Mult_Buf[13].Weight_n = Wgt_0_111;
         Mult_Buf[14].Feature_n = FeatureBuf_112;
         Mult_Buf[14].Weight_n = Wgt_0_112;
         Mult_Buf[15].Feature_n = FeatureBuf_113;
         Mult_Buf[15].Weight_n = Wgt_0_113;
         Mult_Buf[16].Feature_n = FeatureBuf_114;
         Mult_Buf[16].Weight_n = Wgt_0_114;
         Mult_Buf[17].Feature_n = FeatureBuf_115;
         Mult_Buf[17].Weight_n = Wgt_0_115;
         Mult_Buf[18].Feature_n = FeatureBuf_116;
         Mult_Buf[18].Weight_n = Wgt_0_116;
         Mult_Buf[19].Feature_n = FeatureBuf_117;
         Mult_Buf[19].Weight_n = Wgt_0_117;
         Mult_Buf[20].Feature_n = FeatureBuf_118;
         Mult_Buf[20].Weight_n = Wgt_0_118;
         Mult_Buf[21].Feature_n = FeatureBuf_119;
         Mult_Buf[21].Weight_n = Wgt_0_119;
         Mult_Buf[22].Feature_n = FeatureBuf_120;
         Mult_Buf[22].Weight_n = Wgt_0_120;
         Mult_Buf[23].Feature_n = FeatureBuf_121;
         Mult_Buf[23].Weight_n = Wgt_0_121;
         Mult_Buf[24].Feature_n = FeatureBuf_122;
         Mult_Buf[24].Weight_n = Wgt_0_122;
         Mult_Buf[25].Feature_n = FeatureBuf_123;
         Mult_Buf[25].Weight_n = Wgt_0_123;
         Mult_Buf[26].Feature_n = FeatureBuf_124;
         Mult_Buf[26].Weight_n = Wgt_0_124;
         Mult_Buf[27].Feature_n = FeatureBuf_125;
         Mult_Buf[27].Weight_n = Wgt_0_125;
         Mult_Buf[28].Feature_n = FeatureBuf_126;
         Mult_Buf[28].Weight_n = Wgt_0_126;
         Mult_Buf[29].Feature_n = FeatureBuf_127;
         Mult_Buf[29].Weight_n = Wgt_0_127;
         Mult_Buf[30].Feature_n = FeatureBuf_128;
         Mult_Buf[30].Weight_n = Wgt_0_128;
         Mult_Buf[31].Feature_n = FeatureBuf_129;
         Mult_Buf[31].Weight_n = Wgt_0_129;
         Mult_Buf[32].Feature_n = FeatureBuf_130;
         Mult_Buf[32].Weight_n = Wgt_0_130;
         Mult_Buf[33].Feature_n = FeatureBuf_131;
         Mult_Buf[33].Weight_n = Wgt_0_131;
         Mult_Buf[34].Feature_n = FeatureBuf_132;
         Mult_Buf[34].Weight_n = Wgt_0_132;
         Mult_Buf[35].Feature_n = FeatureBuf_133;
         Mult_Buf[35].Weight_n = Wgt_0_133;
         Mult_Buf[36].Feature_n = FeatureBuf_134;
         Mult_Buf[36].Weight_n = Wgt_0_134;
         Mult_Buf[37].Feature_n = FeatureBuf_135;
         Mult_Buf[37].Weight_n = Wgt_0_135;
         Mult_Buf[38].Feature_n = FeatureBuf_136;
         Mult_Buf[38].Weight_n = Wgt_0_136;
         Mult_Buf[39].Feature_n = FeatureBuf_137;
         Mult_Buf[39].Weight_n = Wgt_0_137;
         Mult_Buf[40].Feature_n = FeatureBuf_138;
         Mult_Buf[40].Weight_n = Wgt_0_138;
         Mult_Buf[41].Feature_n = FeatureBuf_139;
         Mult_Buf[41].Weight_n = Wgt_0_139;
         Mult_Buf[42].Feature_n = FeatureBuf_140;
         Mult_Buf[42].Weight_n = Wgt_0_140;
         Mult_Buf[43].Feature_n = FeatureBuf_141;
         Mult_Buf[43].Weight_n = Wgt_0_141;
         Mult_Buf[44].Feature_n = FeatureBuf_142;
         Mult_Buf[44].Weight_n = Wgt_0_142;
         Mult_Buf[45].Feature_n = FeatureBuf_143;
         Mult_Buf[45].Weight_n = Wgt_0_143;
         Mult_Buf[46].Feature_n = FeatureBuf_144;
         Mult_Buf[46].Weight_n = Wgt_0_144;
         Mult_Buf[47].Feature_n = FeatureBuf_145;
         Mult_Buf[47].Weight_n = Wgt_0_145;
         Mult_Buf[48].Feature_n = FeatureBuf_146;
         Mult_Buf[48].Weight_n = Wgt_0_146;
         Mult_Buf[49].Feature_n = FeatureBuf_147;
         Mult_Buf[49].Weight_n = Wgt_0_147;
         Mult_Buf[50].Feature_n = FeatureBuf_148;
         Mult_Buf[50].Weight_n = Wgt_0_148;
         Mult_Buf[51].Feature_n = FeatureBuf_149;
         Mult_Buf[51].Weight_n = Wgt_0_149;
         Mult_Buf[52].Feature_n = FeatureBuf_150;
         Mult_Buf[52].Weight_n = Wgt_0_150;
         Mult_Buf[53].Feature_n = FeatureBuf_151;
         Mult_Buf[53].Weight_n = Wgt_0_151;
         Mult_Buf[54].Feature_n = FeatureBuf_152;
         Mult_Buf[54].Weight_n = Wgt_0_152;
         Mult_Buf[55].Feature_n = FeatureBuf_153;
         Mult_Buf[55].Weight_n = Wgt_0_153;
         Mult_Buf[56].Feature_n = FeatureBuf_154;
         Mult_Buf[56].Weight_n = Wgt_0_154;
         Mult_Buf[57].Feature_n = FeatureBuf_155;
         Mult_Buf[57].Weight_n = Wgt_0_155;
         Mult_Buf[58].Feature_n = FeatureBuf_156;
         Mult_Buf[58].Weight_n = Wgt_0_156;
         Mult_Buf[59].Feature_n = FeatureBuf_157;
         Mult_Buf[59].Weight_n = Wgt_0_157;
         Mult_Buf[60].Feature_n = FeatureBuf_158;
         Mult_Buf[60].Weight_n = Wgt_0_158;
         Mult_Buf[61].Feature_n = FeatureBuf_159;
         Mult_Buf[61].Weight_n = Wgt_0_159;
         Mult_Buf[62].Feature_n = FeatureBuf_160;
         Mult_Buf[62].Weight_n = Wgt_0_160;
         Mult_Buf[63].Feature_n = FeatureBuf_161;
         Mult_Buf[63].Weight_n = Wgt_0_161;
         Mult_Buf[64].Feature_n = FeatureBuf_162;
         Mult_Buf[64].Weight_n = Wgt_0_162;
         Mult_Buf[65].Feature_n = FeatureBuf_163;
         Mult_Buf[65].Weight_n = Wgt_0_163;
         Mult_Buf[66].Feature_n = FeatureBuf_164;
         Mult_Buf[66].Weight_n = Wgt_0_164;
         Mult_Buf[67].Feature_n = FeatureBuf_165;
         Mult_Buf[67].Weight_n = Wgt_0_165;
         Mult_Buf[68].Feature_n = FeatureBuf_166;
         Mult_Buf[68].Weight_n = Wgt_0_166;
         Mult_Buf[69].Feature_n = FeatureBuf_167;
         Mult_Buf[69].Weight_n = Wgt_0_167;
         Mult_Buf[70].Feature_n = FeatureBuf_168;
         Mult_Buf[70].Weight_n = Wgt_0_168;
         Mult_Buf[71].Feature_n = FeatureBuf_169;
         Mult_Buf[71].Weight_n = Wgt_0_169;
         Mult_Buf[72].Feature_n = FeatureBuf_170;
         Mult_Buf[72].Weight_n = Wgt_0_170;
         Mult_Buf[73].Feature_n = FeatureBuf_171;
         Mult_Buf[73].Weight_n = Wgt_0_171;
         Mult_Buf[74].Feature_n = FeatureBuf_172;
         Mult_Buf[74].Weight_n = Wgt_0_172;
         Mult_Buf[75].Feature_n = FeatureBuf_173;
         Mult_Buf[75].Weight_n = Wgt_0_173;
         Mult_Buf[76].Feature_n = FeatureBuf_174;
         Mult_Buf[76].Weight_n = Wgt_0_174;
         Mult_Buf[77].Feature_n = FeatureBuf_175;
         Mult_Buf[77].Weight_n = Wgt_0_175;
         Mult_Buf[78].Feature_n = FeatureBuf_176;
         Mult_Buf[78].Weight_n = Wgt_0_176;
         Mult_Buf[79].Feature_n = FeatureBuf_177;
         Mult_Buf[79].Weight_n = Wgt_0_177;
         Mult_Buf[80].Feature_n = FeatureBuf_178;
         Mult_Buf[80].Weight_n = Wgt_0_178;
         Mult_Buf[81].Feature_n = FeatureBuf_179;
         Mult_Buf[81].Weight_n = Wgt_0_179;
         Mult_Buf[82].Feature_n = FeatureBuf_180;
         Mult_Buf[82].Weight_n = Wgt_0_180;
         Mult_Buf[83].Feature_n = FeatureBuf_181;
         Mult_Buf[83].Weight_n = Wgt_0_181;
         Mult_Buf[84].Feature_n = FeatureBuf_182;
         Mult_Buf[84].Weight_n = Wgt_0_182;
         Mult_Buf[85].Feature_n = FeatureBuf_183;
         Mult_Buf[85].Weight_n = Wgt_0_183;
         Mult_Buf[86].Feature_n = FeatureBuf_184;
         Mult_Buf[86].Weight_n = Wgt_0_184;
         Mult_Buf[87].Feature_n = FeatureBuf_185;
         Mult_Buf[87].Weight_n = Wgt_0_185;
         Mult_Buf[88].Feature_n = FeatureBuf_186;
         Mult_Buf[88].Weight_n = Wgt_0_186;
         Mult_Buf[89].Feature_n = FeatureBuf_187;
         Mult_Buf[89].Weight_n = Wgt_0_187;
         Mult_Buf[90].Feature_n = FeatureBuf_188;
         Mult_Buf[90].Weight_n = Wgt_0_188;
         Mult_Buf[91].Feature_n = FeatureBuf_189;
         Mult_Buf[91].Weight_n = Wgt_0_189;
         Mult_Buf[92].Feature_n = FeatureBuf_190;
         Mult_Buf[92].Weight_n = Wgt_0_190;
         Mult_Buf[93].Feature_n = FeatureBuf_191;
         Mult_Buf[93].Weight_n = Wgt_0_191;
         Mult_Buf[94].Feature_n = FeatureBuf_192;
         Mult_Buf[94].Weight_n = Wgt_0_192;
         Mult_Buf[95].Feature_n = FeatureBuf_193;
         Mult_Buf[95].Weight_n = Wgt_0_193;
         Mult_Buf[96].Feature_n = FeatureBuf_194;
         Mult_Buf[96].Weight_n = Wgt_0_194;
         Mult_Buf[97].Feature_n = FeatureBuf_195;
         Mult_Buf[97].Weight_n = Wgt_0_195;
     end
    4:begin
     nxt_state = 5;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_196;
         Mult_Buf[0].Weight_n = Wgt_0_196;
         Mult_Buf[1].Feature_n = FeatureBuf_197;
         Mult_Buf[1].Weight_n = Wgt_0_197;
         Mult_Buf[2].Feature_n = FeatureBuf_198;
         Mult_Buf[2].Weight_n = Wgt_0_198;
         Mult_Buf[3].Feature_n = FeatureBuf_199;
         Mult_Buf[3].Weight_n = Wgt_0_199;
         Mult_Buf[4].Feature_n = FeatureBuf_200;
         Mult_Buf[4].Weight_n = Wgt_0_200;
         Mult_Buf[5].Feature_n = FeatureBuf_201;
         Mult_Buf[5].Weight_n = Wgt_0_201;
         Mult_Buf[6].Feature_n = FeatureBuf_202;
         Mult_Buf[6].Weight_n = Wgt_0_202;
         Mult_Buf[7].Feature_n = FeatureBuf_203;
         Mult_Buf[7].Weight_n = Wgt_0_203;
         Mult_Buf[8].Feature_n = FeatureBuf_204;
         Mult_Buf[8].Weight_n = Wgt_0_204;
         Mult_Buf[9].Feature_n = FeatureBuf_205;
         Mult_Buf[9].Weight_n = Wgt_0_205;
         Mult_Buf[10].Feature_n = FeatureBuf_206;
         Mult_Buf[10].Weight_n = Wgt_0_206;
         Mult_Buf[11].Feature_n = FeatureBuf_207;
         Mult_Buf[11].Weight_n = Wgt_0_207;
         Mult_Buf[12].Feature_n = FeatureBuf_208;
         Mult_Buf[12].Weight_n = Wgt_0_208;
         Mult_Buf[13].Feature_n = FeatureBuf_209;
         Mult_Buf[13].Weight_n = Wgt_0_209;
         Mult_Buf[14].Feature_n = FeatureBuf_210;
         Mult_Buf[14].Weight_n = Wgt_0_210;
         Mult_Buf[15].Feature_n = FeatureBuf_211;
         Mult_Buf[15].Weight_n = Wgt_0_211;
         Mult_Buf[16].Feature_n = FeatureBuf_212;
         Mult_Buf[16].Weight_n = Wgt_0_212;
         Mult_Buf[17].Feature_n = FeatureBuf_213;
         Mult_Buf[17].Weight_n = Wgt_0_213;
         Mult_Buf[18].Feature_n = FeatureBuf_214;
         Mult_Buf[18].Weight_n = Wgt_0_214;
         Mult_Buf[19].Feature_n = FeatureBuf_215;
         Mult_Buf[19].Weight_n = Wgt_0_215;
         Mult_Buf[20].Feature_n = FeatureBuf_216;
         Mult_Buf[20].Weight_n = Wgt_0_216;
         Mult_Buf[21].Feature_n = FeatureBuf_217;
         Mult_Buf[21].Weight_n = Wgt_0_217;
         Mult_Buf[22].Feature_n = FeatureBuf_218;
         Mult_Buf[22].Weight_n = Wgt_0_218;
         Mult_Buf[23].Feature_n = FeatureBuf_219;
         Mult_Buf[23].Weight_n = Wgt_0_219;
         Mult_Buf[24].Feature_n = FeatureBuf_220;
         Mult_Buf[24].Weight_n = Wgt_0_220;
         Mult_Buf[25].Feature_n = FeatureBuf_221;
         Mult_Buf[25].Weight_n = Wgt_0_221;
         Mult_Buf[26].Feature_n = FeatureBuf_222;
         Mult_Buf[26].Weight_n = Wgt_0_222;
         Mult_Buf[27].Feature_n = FeatureBuf_223;
         Mult_Buf[27].Weight_n = Wgt_0_223;
         Mult_Buf[28].Feature_n = FeatureBuf_224;
         Mult_Buf[28].Weight_n = Wgt_0_224;
         Mult_Buf[29].Feature_n = FeatureBuf_225;
         Mult_Buf[29].Weight_n = Wgt_0_225;
         Mult_Buf[30].Feature_n = FeatureBuf_226;
         Mult_Buf[30].Weight_n = Wgt_0_226;
         Mult_Buf[31].Feature_n = FeatureBuf_227;
         Mult_Buf[31].Weight_n = Wgt_0_227;
         Mult_Buf[32].Feature_n = FeatureBuf_228;
         Mult_Buf[32].Weight_n = Wgt_0_228;
         Mult_Buf[33].Feature_n = FeatureBuf_229;
         Mult_Buf[33].Weight_n = Wgt_0_229;
         Mult_Buf[34].Feature_n = FeatureBuf_230;
         Mult_Buf[34].Weight_n = Wgt_0_230;
         Mult_Buf[35].Feature_n = FeatureBuf_231;
         Mult_Buf[35].Weight_n = Wgt_0_231;
         Mult_Buf[36].Feature_n = FeatureBuf_232;
         Mult_Buf[36].Weight_n = Wgt_0_232;
         Mult_Buf[37].Feature_n = FeatureBuf_233;
         Mult_Buf[37].Weight_n = Wgt_0_233;
         Mult_Buf[38].Feature_n = FeatureBuf_234;
         Mult_Buf[38].Weight_n = Wgt_0_234;
         Mult_Buf[39].Feature_n = FeatureBuf_235;
         Mult_Buf[39].Weight_n = Wgt_0_235;
         Mult_Buf[40].Feature_n = FeatureBuf_236;
         Mult_Buf[40].Weight_n = Wgt_0_236;
         Mult_Buf[41].Feature_n = FeatureBuf_237;
         Mult_Buf[41].Weight_n = Wgt_0_237;
         Mult_Buf[42].Feature_n = FeatureBuf_238;
         Mult_Buf[42].Weight_n = Wgt_0_238;
         Mult_Buf[43].Feature_n = FeatureBuf_239;
         Mult_Buf[43].Weight_n = Wgt_0_239;
         Mult_Buf[44].Feature_n = FeatureBuf_240;
         Mult_Buf[44].Weight_n = Wgt_0_240;
         Mult_Buf[45].Feature_n = FeatureBuf_241;
         Mult_Buf[45].Weight_n = Wgt_0_241;
         Mult_Buf[46].Feature_n = FeatureBuf_242;
         Mult_Buf[46].Weight_n = Wgt_0_242;
         Mult_Buf[47].Feature_n = FeatureBuf_243;
         Mult_Buf[47].Weight_n = Wgt_0_243;
         Mult_Buf[48].Feature_n = FeatureBuf_244;
         Mult_Buf[48].Weight_n = Wgt_0_244;
         Mult_Buf[49].Feature_n = FeatureBuf_245;
         Mult_Buf[49].Weight_n = Wgt_0_245;
         Mult_Buf[50].Feature_n = FeatureBuf_246;
         Mult_Buf[50].Weight_n = Wgt_0_246;
         Mult_Buf[51].Feature_n = FeatureBuf_247;
         Mult_Buf[51].Weight_n = Wgt_0_247;
         Mult_Buf[52].Feature_n = FeatureBuf_248;
         Mult_Buf[52].Weight_n = Wgt_0_248;
         Mult_Buf[53].Feature_n = FeatureBuf_249;
         Mult_Buf[53].Weight_n = Wgt_0_249;
         Mult_Buf[54].Feature_n = FeatureBuf_250;
         Mult_Buf[54].Weight_n = Wgt_0_250;
         Mult_Buf[55].Feature_n = FeatureBuf_251;
         Mult_Buf[55].Weight_n = Wgt_0_251;
         Mult_Buf[56].Feature_n = FeatureBuf_252;
         Mult_Buf[56].Weight_n = Wgt_0_252;
         Mult_Buf[57].Feature_n = FeatureBuf_253;
         Mult_Buf[57].Weight_n = Wgt_0_253;
         Mult_Buf[58].Feature_n = FeatureBuf_254;
         Mult_Buf[58].Weight_n = Wgt_0_254;
         Mult_Buf[59].Feature_n = FeatureBuf_255;
         Mult_Buf[59].Weight_n = Wgt_0_255;
         Mult_Buf[60].Feature_n = FeatureBuf_256;
         Mult_Buf[60].Weight_n = Wgt_0_256;
         Mult_Buf[61].Feature_n = FeatureBuf_257;
         Mult_Buf[61].Weight_n = Wgt_0_257;
         Mult_Buf[62].Feature_n = FeatureBuf_258;
         Mult_Buf[62].Weight_n = Wgt_0_258;
         Mult_Buf[63].Feature_n = FeatureBuf_259;
         Mult_Buf[63].Weight_n = Wgt_0_259;
         Mult_Buf[64].Feature_n = FeatureBuf_260;
         Mult_Buf[64].Weight_n = Wgt_0_260;
         Mult_Buf[65].Feature_n = FeatureBuf_261;
         Mult_Buf[65].Weight_n = Wgt_0_261;
         Mult_Buf[66].Feature_n = FeatureBuf_262;
         Mult_Buf[66].Weight_n = Wgt_0_262;
         Mult_Buf[67].Feature_n = FeatureBuf_263;
         Mult_Buf[67].Weight_n = Wgt_0_263;
         Mult_Buf[68].Feature_n = FeatureBuf_264;
         Mult_Buf[68].Weight_n = Wgt_0_264;
         Mult_Buf[69].Feature_n = FeatureBuf_265;
         Mult_Buf[69].Weight_n = Wgt_0_265;
         Mult_Buf[70].Feature_n = FeatureBuf_266;
         Mult_Buf[70].Weight_n = Wgt_0_266;
         Mult_Buf[71].Feature_n = FeatureBuf_267;
         Mult_Buf[71].Weight_n = Wgt_0_267;
         Mult_Buf[72].Feature_n = FeatureBuf_268;
         Mult_Buf[72].Weight_n = Wgt_0_268;
         Mult_Buf[73].Feature_n = FeatureBuf_269;
         Mult_Buf[73].Weight_n = Wgt_0_269;
         Mult_Buf[74].Feature_n = FeatureBuf_270;
         Mult_Buf[74].Weight_n = Wgt_0_270;
         Mult_Buf[75].Feature_n = FeatureBuf_271;
         Mult_Buf[75].Weight_n = Wgt_0_271;
         Mult_Buf[76].Feature_n = FeatureBuf_272;
         Mult_Buf[76].Weight_n = Wgt_0_272;
         Mult_Buf[77].Feature_n = FeatureBuf_273;
         Mult_Buf[77].Weight_n = Wgt_0_273;
         Mult_Buf[78].Feature_n = FeatureBuf_274;
         Mult_Buf[78].Weight_n = Wgt_0_274;
         Mult_Buf[79].Feature_n = FeatureBuf_275;
         Mult_Buf[79].Weight_n = Wgt_0_275;
         Mult_Buf[80].Feature_n = FeatureBuf_276;
         Mult_Buf[80].Weight_n = Wgt_0_276;
         Mult_Buf[81].Feature_n = FeatureBuf_277;
         Mult_Buf[81].Weight_n = Wgt_0_277;
         Mult_Buf[82].Feature_n = FeatureBuf_278;
         Mult_Buf[82].Weight_n = Wgt_0_278;
         Mult_Buf[83].Feature_n = FeatureBuf_279;
         Mult_Buf[83].Weight_n = Wgt_0_279;
         Mult_Buf[84].Feature_n = FeatureBuf_280;
         Mult_Buf[84].Weight_n = Wgt_0_280;
         Mult_Buf[85].Feature_n = FeatureBuf_281;
         Mult_Buf[85].Weight_n = Wgt_0_281;
         Mult_Buf[86].Feature_n = FeatureBuf_282;
         Mult_Buf[86].Weight_n = Wgt_0_282;
         Mult_Buf[87].Feature_n = FeatureBuf_283;
         Mult_Buf[87].Weight_n = Wgt_0_283;
         Mult_Buf[88].Feature_n = FeatureBuf_284;
         Mult_Buf[88].Weight_n = Wgt_0_284;
         Mult_Buf[89].Feature_n = FeatureBuf_285;
         Mult_Buf[89].Weight_n = Wgt_0_285;
         Mult_Buf[90].Feature_n = FeatureBuf_286;
         Mult_Buf[90].Weight_n = Wgt_0_286;
         Mult_Buf[91].Feature_n = FeatureBuf_287;
         Mult_Buf[91].Weight_n = Wgt_0_287;
         Mult_Buf[92].Feature_n = FeatureBuf_288;
         Mult_Buf[92].Weight_n = Wgt_0_288;
         Mult_Buf[93].Feature_n = FeatureBuf_289;
         Mult_Buf[93].Weight_n = Wgt_0_289;
         Mult_Buf[94].Feature_n = FeatureBuf_290;
         Mult_Buf[94].Weight_n = Wgt_0_290;
         Mult_Buf[95].Feature_n = FeatureBuf_291;
         Mult_Buf[95].Weight_n = Wgt_0_291;
         Mult_Buf[96].Feature_n = FeatureBuf_292;
         Mult_Buf[96].Weight_n = Wgt_0_292;
         Mult_Buf[97].Feature_n = FeatureBuf_293;
         Mult_Buf[97].Weight_n = Wgt_0_293;
     end
    5:begin
     nxt_state = 6;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_294;
         Mult_Buf[0].Weight_n = Wgt_0_294;
         Mult_Buf[1].Feature_n = FeatureBuf_295;
         Mult_Buf[1].Weight_n = Wgt_0_295;
         Mult_Buf[2].Feature_n = FeatureBuf_296;
         Mult_Buf[2].Weight_n = Wgt_0_296;
         Mult_Buf[3].Feature_n = FeatureBuf_297;
         Mult_Buf[3].Weight_n = Wgt_0_297;
         Mult_Buf[4].Feature_n = FeatureBuf_298;
         Mult_Buf[4].Weight_n = Wgt_0_298;
         Mult_Buf[5].Feature_n = FeatureBuf_299;
         Mult_Buf[5].Weight_n = Wgt_0_299;
         Mult_Buf[6].Feature_n = FeatureBuf_300;
         Mult_Buf[6].Weight_n = Wgt_0_300;
         Mult_Buf[7].Feature_n = FeatureBuf_301;
         Mult_Buf[7].Weight_n = Wgt_0_301;
         Mult_Buf[8].Feature_n = FeatureBuf_302;
         Mult_Buf[8].Weight_n = Wgt_0_302;
         Mult_Buf[9].Feature_n = FeatureBuf_303;
         Mult_Buf[9].Weight_n = Wgt_0_303;
         Mult_Buf[10].Feature_n = FeatureBuf_304;
         Mult_Buf[10].Weight_n = Wgt_0_304;
         Mult_Buf[11].Feature_n = FeatureBuf_305;
         Mult_Buf[11].Weight_n = Wgt_0_305;
         Mult_Buf[12].Feature_n = FeatureBuf_306;
         Mult_Buf[12].Weight_n = Wgt_0_306;
         Mult_Buf[13].Feature_n = FeatureBuf_307;
         Mult_Buf[13].Weight_n = Wgt_0_307;
         Mult_Buf[14].Feature_n = FeatureBuf_308;
         Mult_Buf[14].Weight_n = Wgt_0_308;
         Mult_Buf[15].Feature_n = FeatureBuf_309;
         Mult_Buf[15].Weight_n = Wgt_0_309;
         Mult_Buf[16].Feature_n = FeatureBuf_310;
         Mult_Buf[16].Weight_n = Wgt_0_310;
         Mult_Buf[17].Feature_n = FeatureBuf_311;
         Mult_Buf[17].Weight_n = Wgt_0_311;
         Mult_Buf[18].Feature_n = FeatureBuf_312;
         Mult_Buf[18].Weight_n = Wgt_0_312;
         Mult_Buf[19].Feature_n = FeatureBuf_313;
         Mult_Buf[19].Weight_n = Wgt_0_313;
         Mult_Buf[20].Feature_n = FeatureBuf_314;
         Mult_Buf[20].Weight_n = Wgt_0_314;
         Mult_Buf[21].Feature_n = FeatureBuf_315;
         Mult_Buf[21].Weight_n = Wgt_0_315;
         Mult_Buf[22].Feature_n = FeatureBuf_316;
         Mult_Buf[22].Weight_n = Wgt_0_316;
         Mult_Buf[23].Feature_n = FeatureBuf_317;
         Mult_Buf[23].Weight_n = Wgt_0_317;
         Mult_Buf[24].Feature_n = FeatureBuf_318;
         Mult_Buf[24].Weight_n = Wgt_0_318;
         Mult_Buf[25].Feature_n = FeatureBuf_319;
         Mult_Buf[25].Weight_n = Wgt_0_319;
         Mult_Buf[26].Feature_n = FeatureBuf_320;
         Mult_Buf[26].Weight_n = Wgt_0_320;
         Mult_Buf[27].Feature_n = FeatureBuf_321;
         Mult_Buf[27].Weight_n = Wgt_0_321;
         Mult_Buf[28].Feature_n = FeatureBuf_322;
         Mult_Buf[28].Weight_n = Wgt_0_322;
         Mult_Buf[29].Feature_n = FeatureBuf_323;
         Mult_Buf[29].Weight_n = Wgt_0_323;
         Mult_Buf[30].Feature_n = FeatureBuf_324;
         Mult_Buf[30].Weight_n = Wgt_0_324;
         Mult_Buf[31].Feature_n = FeatureBuf_325;
         Mult_Buf[31].Weight_n = Wgt_0_325;
         Mult_Buf[32].Feature_n = FeatureBuf_326;
         Mult_Buf[32].Weight_n = Wgt_0_326;
         Mult_Buf[33].Feature_n = FeatureBuf_327;
         Mult_Buf[33].Weight_n = Wgt_0_327;
         Mult_Buf[34].Feature_n = FeatureBuf_328;
         Mult_Buf[34].Weight_n = Wgt_0_328;
         Mult_Buf[35].Feature_n = FeatureBuf_329;
         Mult_Buf[35].Weight_n = Wgt_0_329;
         Mult_Buf[36].Feature_n = FeatureBuf_330;
         Mult_Buf[36].Weight_n = Wgt_0_330;
         Mult_Buf[37].Feature_n = FeatureBuf_331;
         Mult_Buf[37].Weight_n = Wgt_0_331;
         Mult_Buf[38].Feature_n = FeatureBuf_332;
         Mult_Buf[38].Weight_n = Wgt_0_332;
         Mult_Buf[39].Feature_n = FeatureBuf_333;
         Mult_Buf[39].Weight_n = Wgt_0_333;
         Mult_Buf[40].Feature_n = FeatureBuf_334;
         Mult_Buf[40].Weight_n = Wgt_0_334;
         Mult_Buf[41].Feature_n = FeatureBuf_335;
         Mult_Buf[41].Weight_n = Wgt_0_335;
         Mult_Buf[42].Feature_n = FeatureBuf_336;
         Mult_Buf[42].Weight_n = Wgt_0_336;
         Mult_Buf[43].Feature_n = FeatureBuf_337;
         Mult_Buf[43].Weight_n = Wgt_0_337;
         Mult_Buf[44].Feature_n = FeatureBuf_338;
         Mult_Buf[44].Weight_n = Wgt_0_338;
         Mult_Buf[45].Feature_n = FeatureBuf_339;
         Mult_Buf[45].Weight_n = Wgt_0_339;
         Mult_Buf[46].Feature_n = FeatureBuf_340;
         Mult_Buf[46].Weight_n = Wgt_0_340;
         Mult_Buf[47].Feature_n = FeatureBuf_341;
         Mult_Buf[47].Weight_n = Wgt_0_341;
         Mult_Buf[48].Feature_n = FeatureBuf_342;
         Mult_Buf[48].Weight_n = Wgt_0_342;
         Mult_Buf[49].Feature_n = FeatureBuf_343;
         Mult_Buf[49].Weight_n = Wgt_0_343;
         Mult_Buf[50].Feature_n = FeatureBuf_344;
         Mult_Buf[50].Weight_n = Wgt_0_344;
         Mult_Buf[51].Feature_n = FeatureBuf_345;
         Mult_Buf[51].Weight_n = Wgt_0_345;
         Mult_Buf[52].Feature_n = FeatureBuf_346;
         Mult_Buf[52].Weight_n = Wgt_0_346;
         Mult_Buf[53].Feature_n = FeatureBuf_347;
         Mult_Buf[53].Weight_n = Wgt_0_347;
         Mult_Buf[54].Feature_n = FeatureBuf_348;
         Mult_Buf[54].Weight_n = Wgt_0_348;
         Mult_Buf[55].Feature_n = FeatureBuf_349;
         Mult_Buf[55].Weight_n = Wgt_0_349;
         Mult_Buf[56].Feature_n = FeatureBuf_350;
         Mult_Buf[56].Weight_n = Wgt_0_350;
         Mult_Buf[57].Feature_n = FeatureBuf_351;
         Mult_Buf[57].Weight_n = Wgt_0_351;
         Mult_Buf[58].Feature_n = FeatureBuf_352;
         Mult_Buf[58].Weight_n = Wgt_0_352;
         Mult_Buf[59].Feature_n = FeatureBuf_353;
         Mult_Buf[59].Weight_n = Wgt_0_353;
         Mult_Buf[60].Feature_n = FeatureBuf_354;
         Mult_Buf[60].Weight_n = Wgt_0_354;
         Mult_Buf[61].Feature_n = FeatureBuf_355;
         Mult_Buf[61].Weight_n = Wgt_0_355;
         Mult_Buf[62].Feature_n = FeatureBuf_356;
         Mult_Buf[62].Weight_n = Wgt_0_356;
         Mult_Buf[63].Feature_n = FeatureBuf_357;
         Mult_Buf[63].Weight_n = Wgt_0_357;
         Mult_Buf[64].Feature_n = FeatureBuf_358;
         Mult_Buf[64].Weight_n = Wgt_0_358;
         Mult_Buf[65].Feature_n = FeatureBuf_359;
         Mult_Buf[65].Weight_n = Wgt_0_359;
         Mult_Buf[66].Feature_n = FeatureBuf_360;
         Mult_Buf[66].Weight_n = Wgt_0_360;
         Mult_Buf[67].Feature_n = FeatureBuf_361;
         Mult_Buf[67].Weight_n = Wgt_0_361;
         Mult_Buf[68].Feature_n = FeatureBuf_362;
         Mult_Buf[68].Weight_n = Wgt_0_362;
         Mult_Buf[69].Feature_n = FeatureBuf_363;
         Mult_Buf[69].Weight_n = Wgt_0_363;
         Mult_Buf[70].Feature_n = FeatureBuf_364;
         Mult_Buf[70].Weight_n = Wgt_0_364;
         Mult_Buf[71].Feature_n = FeatureBuf_365;
         Mult_Buf[71].Weight_n = Wgt_0_365;
         Mult_Buf[72].Feature_n = FeatureBuf_366;
         Mult_Buf[72].Weight_n = Wgt_0_366;
         Mult_Buf[73].Feature_n = FeatureBuf_367;
         Mult_Buf[73].Weight_n = Wgt_0_367;
         Mult_Buf[74].Feature_n = FeatureBuf_368;
         Mult_Buf[74].Weight_n = Wgt_0_368;
         Mult_Buf[75].Feature_n = FeatureBuf_369;
         Mult_Buf[75].Weight_n = Wgt_0_369;
         Mult_Buf[76].Feature_n = FeatureBuf_370;
         Mult_Buf[76].Weight_n = Wgt_0_370;
         Mult_Buf[77].Feature_n = FeatureBuf_371;
         Mult_Buf[77].Weight_n = Wgt_0_371;
         Mult_Buf[78].Feature_n = FeatureBuf_372;
         Mult_Buf[78].Weight_n = Wgt_0_372;
         Mult_Buf[79].Feature_n = FeatureBuf_373;
         Mult_Buf[79].Weight_n = Wgt_0_373;
         Mult_Buf[80].Feature_n = FeatureBuf_374;
         Mult_Buf[80].Weight_n = Wgt_0_374;
         Mult_Buf[81].Feature_n = FeatureBuf_375;
         Mult_Buf[81].Weight_n = Wgt_0_375;
         Mult_Buf[82].Feature_n = FeatureBuf_376;
         Mult_Buf[82].Weight_n = Wgt_0_376;
         Mult_Buf[83].Feature_n = FeatureBuf_377;
         Mult_Buf[83].Weight_n = Wgt_0_377;
         Mult_Buf[84].Feature_n = FeatureBuf_378;
         Mult_Buf[84].Weight_n = Wgt_0_378;
         Mult_Buf[85].Feature_n = FeatureBuf_379;
         Mult_Buf[85].Weight_n = Wgt_0_379;
         Mult_Buf[86].Feature_n = FeatureBuf_380;
         Mult_Buf[86].Weight_n = Wgt_0_380;
         Mult_Buf[87].Feature_n = FeatureBuf_381;
         Mult_Buf[87].Weight_n = Wgt_0_381;
         Mult_Buf[88].Feature_n = FeatureBuf_382;
         Mult_Buf[88].Weight_n = Wgt_0_382;
         Mult_Buf[89].Feature_n = FeatureBuf_383;
         Mult_Buf[89].Weight_n = Wgt_0_383;
         Mult_Buf[90].Feature_n = FeatureBuf_384;
         Mult_Buf[90].Weight_n = Wgt_0_384;
         Mult_Buf[91].Feature_n = FeatureBuf_385;
         Mult_Buf[91].Weight_n = Wgt_0_385;
         Mult_Buf[92].Feature_n = FeatureBuf_386;
         Mult_Buf[92].Weight_n = Wgt_0_386;
         Mult_Buf[93].Feature_n = FeatureBuf_387;
         Mult_Buf[93].Weight_n = Wgt_0_387;
         Mult_Buf[94].Feature_n = FeatureBuf_388;
         Mult_Buf[94].Weight_n = Wgt_0_388;
         Mult_Buf[95].Feature_n = FeatureBuf_389;
         Mult_Buf[95].Weight_n = Wgt_0_389;
         Mult_Buf[96].Feature_n = FeatureBuf_390;
         Mult_Buf[96].Weight_n = Wgt_0_390;
         Mult_Buf[97].Feature_n = FeatureBuf_391;
         Mult_Buf[97].Weight_n = Wgt_0_391;
     end
    6:begin
     nxt_state = 7;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_392;
         Mult_Buf[0].Weight_n = Wgt_0_392;
         Mult_Buf[1].Feature_n = FeatureBuf_393;
         Mult_Buf[1].Weight_n = Wgt_0_393;
         Mult_Buf[2].Feature_n = FeatureBuf_394;
         Mult_Buf[2].Weight_n = Wgt_0_394;
         Mult_Buf[3].Feature_n = FeatureBuf_395;
         Mult_Buf[3].Weight_n = Wgt_0_395;
         Mult_Buf[4].Feature_n = FeatureBuf_396;
         Mult_Buf[4].Weight_n = Wgt_0_396;
         Mult_Buf[5].Feature_n = FeatureBuf_397;
         Mult_Buf[5].Weight_n = Wgt_0_397;
         Mult_Buf[6].Feature_n = FeatureBuf_398;
         Mult_Buf[6].Weight_n = Wgt_0_398;
         Mult_Buf[7].Feature_n = FeatureBuf_399;
         Mult_Buf[7].Weight_n = Wgt_0_399;
         Mult_Buf[8].Feature_n = FeatureBuf_400;
         Mult_Buf[8].Weight_n = Wgt_0_400;
         Mult_Buf[9].Feature_n = FeatureBuf_401;
         Mult_Buf[9].Weight_n = Wgt_0_401;
         Mult_Buf[10].Feature_n = FeatureBuf_402;
         Mult_Buf[10].Weight_n = Wgt_0_402;
         Mult_Buf[11].Feature_n = FeatureBuf_403;
         Mult_Buf[11].Weight_n = Wgt_0_403;
         Mult_Buf[12].Feature_n = FeatureBuf_404;
         Mult_Buf[12].Weight_n = Wgt_0_404;
         Mult_Buf[13].Feature_n = FeatureBuf_405;
         Mult_Buf[13].Weight_n = Wgt_0_405;
         Mult_Buf[14].Feature_n = FeatureBuf_406;
         Mult_Buf[14].Weight_n = Wgt_0_406;
         Mult_Buf[15].Feature_n = FeatureBuf_407;
         Mult_Buf[15].Weight_n = Wgt_0_407;
         Mult_Buf[16].Feature_n = FeatureBuf_408;
         Mult_Buf[16].Weight_n = Wgt_0_408;
         Mult_Buf[17].Feature_n = FeatureBuf_409;
         Mult_Buf[17].Weight_n = Wgt_0_409;
         Mult_Buf[18].Feature_n = FeatureBuf_410;
         Mult_Buf[18].Weight_n = Wgt_0_410;
         Mult_Buf[19].Feature_n = FeatureBuf_411;
         Mult_Buf[19].Weight_n = Wgt_0_411;
         Mult_Buf[20].Feature_n = FeatureBuf_412;
         Mult_Buf[20].Weight_n = Wgt_0_412;
         Mult_Buf[21].Feature_n = FeatureBuf_413;
         Mult_Buf[21].Weight_n = Wgt_0_413;
         Mult_Buf[22].Feature_n = FeatureBuf_414;
         Mult_Buf[22].Weight_n = Wgt_0_414;
         Mult_Buf[23].Feature_n = FeatureBuf_415;
         Mult_Buf[23].Weight_n = Wgt_0_415;
         Mult_Buf[24].Feature_n = FeatureBuf_416;
         Mult_Buf[24].Weight_n = Wgt_0_416;
         Mult_Buf[25].Feature_n = FeatureBuf_417;
         Mult_Buf[25].Weight_n = Wgt_0_417;
         Mult_Buf[26].Feature_n = FeatureBuf_418;
         Mult_Buf[26].Weight_n = Wgt_0_418;
         Mult_Buf[27].Feature_n = FeatureBuf_419;
         Mult_Buf[27].Weight_n = Wgt_0_419;
         Mult_Buf[28].Feature_n = FeatureBuf_420;
         Mult_Buf[28].Weight_n = Wgt_0_420;
         Mult_Buf[29].Feature_n = FeatureBuf_421;
         Mult_Buf[29].Weight_n = Wgt_0_421;
         Mult_Buf[30].Feature_n = FeatureBuf_422;
         Mult_Buf[30].Weight_n = Wgt_0_422;
         Mult_Buf[31].Feature_n = FeatureBuf_423;
         Mult_Buf[31].Weight_n = Wgt_0_423;
         Mult_Buf[32].Feature_n = FeatureBuf_424;
         Mult_Buf[32].Weight_n = Wgt_0_424;
         Mult_Buf[33].Feature_n = FeatureBuf_425;
         Mult_Buf[33].Weight_n = Wgt_0_425;
         Mult_Buf[34].Feature_n = FeatureBuf_426;
         Mult_Buf[34].Weight_n = Wgt_0_426;
         Mult_Buf[35].Feature_n = FeatureBuf_427;
         Mult_Buf[35].Weight_n = Wgt_0_427;
         Mult_Buf[36].Feature_n = FeatureBuf_428;
         Mult_Buf[36].Weight_n = Wgt_0_428;
         Mult_Buf[37].Feature_n = FeatureBuf_429;
         Mult_Buf[37].Weight_n = Wgt_0_429;
         Mult_Buf[38].Feature_n = FeatureBuf_430;
         Mult_Buf[38].Weight_n = Wgt_0_430;
         Mult_Buf[39].Feature_n = FeatureBuf_431;
         Mult_Buf[39].Weight_n = Wgt_0_431;
         Mult_Buf[40].Feature_n = FeatureBuf_432;
         Mult_Buf[40].Weight_n = Wgt_0_432;
         Mult_Buf[41].Feature_n = FeatureBuf_433;
         Mult_Buf[41].Weight_n = Wgt_0_433;
         Mult_Buf[42].Feature_n = FeatureBuf_434;
         Mult_Buf[42].Weight_n = Wgt_0_434;
         Mult_Buf[43].Feature_n = FeatureBuf_435;
         Mult_Buf[43].Weight_n = Wgt_0_435;
         Mult_Buf[44].Feature_n = FeatureBuf_436;
         Mult_Buf[44].Weight_n = Wgt_0_436;
         Mult_Buf[45].Feature_n = FeatureBuf_437;
         Mult_Buf[45].Weight_n = Wgt_0_437;
         Mult_Buf[46].Feature_n = FeatureBuf_438;
         Mult_Buf[46].Weight_n = Wgt_0_438;
         Mult_Buf[47].Feature_n = FeatureBuf_439;
         Mult_Buf[47].Weight_n = Wgt_0_439;
         Mult_Buf[48].Feature_n = FeatureBuf_440;
         Mult_Buf[48].Weight_n = Wgt_0_440;
         Mult_Buf[49].Feature_n = FeatureBuf_441;
         Mult_Buf[49].Weight_n = Wgt_0_441;
         Mult_Buf[50].Feature_n = FeatureBuf_442;
         Mult_Buf[50].Weight_n = Wgt_0_442;
         Mult_Buf[51].Feature_n = FeatureBuf_443;
         Mult_Buf[51].Weight_n = Wgt_0_443;
         Mult_Buf[52].Feature_n = FeatureBuf_444;
         Mult_Buf[52].Weight_n = Wgt_0_444;
         Mult_Buf[53].Feature_n = FeatureBuf_445;
         Mult_Buf[53].Weight_n = Wgt_0_445;
         Mult_Buf[54].Feature_n = FeatureBuf_446;
         Mult_Buf[54].Weight_n = Wgt_0_446;
         Mult_Buf[55].Feature_n = FeatureBuf_447;
         Mult_Buf[55].Weight_n = Wgt_0_447;
         Mult_Buf[56].Feature_n = FeatureBuf_448;
         Mult_Buf[56].Weight_n = Wgt_0_448;
         Mult_Buf[57].Feature_n = FeatureBuf_449;
         Mult_Buf[57].Weight_n = Wgt_0_449;
         Mult_Buf[58].Feature_n = FeatureBuf_450;
         Mult_Buf[58].Weight_n = Wgt_0_450;
         Mult_Buf[59].Feature_n = FeatureBuf_451;
         Mult_Buf[59].Weight_n = Wgt_0_451;
         Mult_Buf[60].Feature_n = FeatureBuf_452;
         Mult_Buf[60].Weight_n = Wgt_0_452;
         Mult_Buf[61].Feature_n = FeatureBuf_453;
         Mult_Buf[61].Weight_n = Wgt_0_453;
         Mult_Buf[62].Feature_n = FeatureBuf_454;
         Mult_Buf[62].Weight_n = Wgt_0_454;
         Mult_Buf[63].Feature_n = FeatureBuf_455;
         Mult_Buf[63].Weight_n = Wgt_0_455;
         Mult_Buf[64].Feature_n = FeatureBuf_456;
         Mult_Buf[64].Weight_n = Wgt_0_456;
         Mult_Buf[65].Feature_n = FeatureBuf_457;
         Mult_Buf[65].Weight_n = Wgt_0_457;
         Mult_Buf[66].Feature_n = FeatureBuf_458;
         Mult_Buf[66].Weight_n = Wgt_0_458;
         Mult_Buf[67].Feature_n = FeatureBuf_459;
         Mult_Buf[67].Weight_n = Wgt_0_459;
         Mult_Buf[68].Feature_n = FeatureBuf_460;
         Mult_Buf[68].Weight_n = Wgt_0_460;
         Mult_Buf[69].Feature_n = FeatureBuf_461;
         Mult_Buf[69].Weight_n = Wgt_0_461;
         Mult_Buf[70].Feature_n = FeatureBuf_462;
         Mult_Buf[70].Weight_n = Wgt_0_462;
         Mult_Buf[71].Feature_n = FeatureBuf_463;
         Mult_Buf[71].Weight_n = Wgt_0_463;
         Mult_Buf[72].Feature_n = FeatureBuf_464;
         Mult_Buf[72].Weight_n = Wgt_0_464;
         Mult_Buf[73].Feature_n = FeatureBuf_465;
         Mult_Buf[73].Weight_n = Wgt_0_465;
         Mult_Buf[74].Feature_n = FeatureBuf_466;
         Mult_Buf[74].Weight_n = Wgt_0_466;
         Mult_Buf[75].Feature_n = FeatureBuf_467;
         Mult_Buf[75].Weight_n = Wgt_0_467;
         Mult_Buf[76].Feature_n = FeatureBuf_468;
         Mult_Buf[76].Weight_n = Wgt_0_468;
         Mult_Buf[77].Feature_n = FeatureBuf_469;
         Mult_Buf[77].Weight_n = Wgt_0_469;
         Mult_Buf[78].Feature_n = FeatureBuf_470;
         Mult_Buf[78].Weight_n = Wgt_0_470;
         Mult_Buf[79].Feature_n = FeatureBuf_471;
         Mult_Buf[79].Weight_n = Wgt_0_471;
         Mult_Buf[80].Feature_n = FeatureBuf_472;
         Mult_Buf[80].Weight_n = Wgt_0_472;
         Mult_Buf[81].Feature_n = FeatureBuf_473;
         Mult_Buf[81].Weight_n = Wgt_0_473;
         Mult_Buf[82].Feature_n = FeatureBuf_474;
         Mult_Buf[82].Weight_n = Wgt_0_474;
         Mult_Buf[83].Feature_n = FeatureBuf_475;
         Mult_Buf[83].Weight_n = Wgt_0_475;
         Mult_Buf[84].Feature_n = FeatureBuf_476;
         Mult_Buf[84].Weight_n = Wgt_0_476;
         Mult_Buf[85].Feature_n = FeatureBuf_477;
         Mult_Buf[85].Weight_n = Wgt_0_477;
         Mult_Buf[86].Feature_n = FeatureBuf_478;
         Mult_Buf[86].Weight_n = Wgt_0_478;
         Mult_Buf[87].Feature_n = FeatureBuf_479;
         Mult_Buf[87].Weight_n = Wgt_0_479;
         Mult_Buf[88].Feature_n = FeatureBuf_480;
         Mult_Buf[88].Weight_n = Wgt_0_480;
         Mult_Buf[89].Feature_n = FeatureBuf_481;
         Mult_Buf[89].Weight_n = Wgt_0_481;
         Mult_Buf[90].Feature_n = FeatureBuf_482;
         Mult_Buf[90].Weight_n = Wgt_0_482;
         Mult_Buf[91].Feature_n = FeatureBuf_483;
         Mult_Buf[91].Weight_n = Wgt_0_483;
         Mult_Buf[92].Feature_n = FeatureBuf_484;
         Mult_Buf[92].Weight_n = Wgt_0_484;
         Mult_Buf[93].Feature_n = FeatureBuf_485;
         Mult_Buf[93].Weight_n = Wgt_0_485;
         Mult_Buf[94].Feature_n = FeatureBuf_486;
         Mult_Buf[94].Weight_n = Wgt_0_486;
         Mult_Buf[95].Feature_n = FeatureBuf_487;
         Mult_Buf[95].Weight_n = Wgt_0_487;
         Mult_Buf[96].Feature_n = FeatureBuf_488;
         Mult_Buf[96].Weight_n = Wgt_0_488;
         Mult_Buf[97].Feature_n = FeatureBuf_489;
         Mult_Buf[97].Weight_n = Wgt_0_489;
     end
    7:begin
     nxt_state = 8;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_490;
         Mult_Buf[0].Weight_n = Wgt_0_490;
         Mult_Buf[1].Feature_n = FeatureBuf_491;
         Mult_Buf[1].Weight_n = Wgt_0_491;
         Mult_Buf[2].Feature_n = FeatureBuf_492;
         Mult_Buf[2].Weight_n = Wgt_0_492;
         Mult_Buf[3].Feature_n = FeatureBuf_493;
         Mult_Buf[3].Weight_n = Wgt_0_493;
         Mult_Buf[4].Feature_n = FeatureBuf_494;
         Mult_Buf[4].Weight_n = Wgt_0_494;
         Mult_Buf[5].Feature_n = FeatureBuf_495;
         Mult_Buf[5].Weight_n = Wgt_0_495;
         Mult_Buf[6].Feature_n = FeatureBuf_496;
         Mult_Buf[6].Weight_n = Wgt_0_496;
         Mult_Buf[7].Feature_n = FeatureBuf_497;
         Mult_Buf[7].Weight_n = Wgt_0_497;
         Mult_Buf[8].Feature_n = FeatureBuf_498;
         Mult_Buf[8].Weight_n = Wgt_0_498;
         Mult_Buf[9].Feature_n = FeatureBuf_499;
         Mult_Buf[9].Weight_n = Wgt_0_499;
         Mult_Buf[10].Feature_n = FeatureBuf_500;
         Mult_Buf[10].Weight_n = Wgt_0_500;
         Mult_Buf[11].Feature_n = FeatureBuf_501;
         Mult_Buf[11].Weight_n = Wgt_0_501;
         Mult_Buf[12].Feature_n = FeatureBuf_502;
         Mult_Buf[12].Weight_n = Wgt_0_502;
         Mult_Buf[13].Feature_n = FeatureBuf_503;
         Mult_Buf[13].Weight_n = Wgt_0_503;
         Mult_Buf[14].Feature_n = FeatureBuf_504;
         Mult_Buf[14].Weight_n = Wgt_0_504;
         Mult_Buf[15].Feature_n = FeatureBuf_505;
         Mult_Buf[15].Weight_n = Wgt_0_505;
         Mult_Buf[16].Feature_n = FeatureBuf_506;
         Mult_Buf[16].Weight_n = Wgt_0_506;
         Mult_Buf[17].Feature_n = FeatureBuf_507;
         Mult_Buf[17].Weight_n = Wgt_0_507;
         Mult_Buf[18].Feature_n = FeatureBuf_508;
         Mult_Buf[18].Weight_n = Wgt_0_508;
         Mult_Buf[19].Feature_n = FeatureBuf_509;
         Mult_Buf[19].Weight_n = Wgt_0_509;
         Mult_Buf[20].Feature_n = FeatureBuf_510;
         Mult_Buf[20].Weight_n = Wgt_0_510;
         Mult_Buf[21].Feature_n = FeatureBuf_511;
         Mult_Buf[21].Weight_n = Wgt_0_511;
         Mult_Buf[22].Feature_n = FeatureBuf_512;
         Mult_Buf[22].Weight_n = Wgt_0_512;
         Mult_Buf[23].Feature_n = FeatureBuf_513;
         Mult_Buf[23].Weight_n = Wgt_0_513;
         Mult_Buf[24].Feature_n = FeatureBuf_514;
         Mult_Buf[24].Weight_n = Wgt_0_514;
         Mult_Buf[25].Feature_n = FeatureBuf_515;
         Mult_Buf[25].Weight_n = Wgt_0_515;
         Mult_Buf[26].Feature_n = FeatureBuf_516;
         Mult_Buf[26].Weight_n = Wgt_0_516;
         Mult_Buf[27].Feature_n = FeatureBuf_517;
         Mult_Buf[27].Weight_n = Wgt_0_517;
         Mult_Buf[28].Feature_n = FeatureBuf_518;
         Mult_Buf[28].Weight_n = Wgt_0_518;
         Mult_Buf[29].Feature_n = FeatureBuf_519;
         Mult_Buf[29].Weight_n = Wgt_0_519;
         Mult_Buf[30].Feature_n = FeatureBuf_520;
         Mult_Buf[30].Weight_n = Wgt_0_520;
         Mult_Buf[31].Feature_n = FeatureBuf_521;
         Mult_Buf[31].Weight_n = Wgt_0_521;
         Mult_Buf[32].Feature_n = FeatureBuf_522;
         Mult_Buf[32].Weight_n = Wgt_0_522;
         Mult_Buf[33].Feature_n = FeatureBuf_523;
         Mult_Buf[33].Weight_n = Wgt_0_523;
         Mult_Buf[34].Feature_n = FeatureBuf_524;
         Mult_Buf[34].Weight_n = Wgt_0_524;
         Mult_Buf[35].Feature_n = FeatureBuf_525;
         Mult_Buf[35].Weight_n = Wgt_0_525;
         Mult_Buf[36].Feature_n = FeatureBuf_526;
         Mult_Buf[36].Weight_n = Wgt_0_526;
         Mult_Buf[37].Feature_n = FeatureBuf_527;
         Mult_Buf[37].Weight_n = Wgt_0_527;
         Mult_Buf[38].Feature_n = FeatureBuf_528;
         Mult_Buf[38].Weight_n = Wgt_0_528;
         Mult_Buf[39].Feature_n = FeatureBuf_529;
         Mult_Buf[39].Weight_n = Wgt_0_529;
         Mult_Buf[40].Feature_n = FeatureBuf_530;
         Mult_Buf[40].Weight_n = Wgt_0_530;
         Mult_Buf[41].Feature_n = FeatureBuf_531;
         Mult_Buf[41].Weight_n = Wgt_0_531;
         Mult_Buf[42].Feature_n = FeatureBuf_532;
         Mult_Buf[42].Weight_n = Wgt_0_532;
         Mult_Buf[43].Feature_n = FeatureBuf_533;
         Mult_Buf[43].Weight_n = Wgt_0_533;
         Mult_Buf[44].Feature_n = FeatureBuf_534;
         Mult_Buf[44].Weight_n = Wgt_0_534;
         Mult_Buf[45].Feature_n = FeatureBuf_535;
         Mult_Buf[45].Weight_n = Wgt_0_535;
         Mult_Buf[46].Feature_n = FeatureBuf_536;
         Mult_Buf[46].Weight_n = Wgt_0_536;
         Mult_Buf[47].Feature_n = FeatureBuf_537;
         Mult_Buf[47].Weight_n = Wgt_0_537;
         Mult_Buf[48].Feature_n = FeatureBuf_538;
         Mult_Buf[48].Weight_n = Wgt_0_538;
         Mult_Buf[49].Feature_n = FeatureBuf_539;
         Mult_Buf[49].Weight_n = Wgt_0_539;
         Mult_Buf[50].Feature_n = FeatureBuf_540;
         Mult_Buf[50].Weight_n = Wgt_0_540;
         Mult_Buf[51].Feature_n = FeatureBuf_541;
         Mult_Buf[51].Weight_n = Wgt_0_541;
         Mult_Buf[52].Feature_n = FeatureBuf_542;
         Mult_Buf[52].Weight_n = Wgt_0_542;
         Mult_Buf[53].Feature_n = FeatureBuf_543;
         Mult_Buf[53].Weight_n = Wgt_0_543;
         Mult_Buf[54].Feature_n = FeatureBuf_544;
         Mult_Buf[54].Weight_n = Wgt_0_544;
         Mult_Buf[55].Feature_n = FeatureBuf_545;
         Mult_Buf[55].Weight_n = Wgt_0_545;
         Mult_Buf[56].Feature_n = FeatureBuf_546;
         Mult_Buf[56].Weight_n = Wgt_0_546;
         Mult_Buf[57].Feature_n = FeatureBuf_547;
         Mult_Buf[57].Weight_n = Wgt_0_547;
         Mult_Buf[58].Feature_n = FeatureBuf_548;
         Mult_Buf[58].Weight_n = Wgt_0_548;
         Mult_Buf[59].Feature_n = FeatureBuf_549;
         Mult_Buf[59].Weight_n = Wgt_0_549;
         Mult_Buf[60].Feature_n = FeatureBuf_550;
         Mult_Buf[60].Weight_n = Wgt_0_550;
         Mult_Buf[61].Feature_n = FeatureBuf_551;
         Mult_Buf[61].Weight_n = Wgt_0_551;
         Mult_Buf[62].Feature_n = FeatureBuf_552;
         Mult_Buf[62].Weight_n = Wgt_0_552;
         Mult_Buf[63].Feature_n = FeatureBuf_553;
         Mult_Buf[63].Weight_n = Wgt_0_553;
         Mult_Buf[64].Feature_n = FeatureBuf_554;
         Mult_Buf[64].Weight_n = Wgt_0_554;
         Mult_Buf[65].Feature_n = FeatureBuf_555;
         Mult_Buf[65].Weight_n = Wgt_0_555;
         Mult_Buf[66].Feature_n = FeatureBuf_556;
         Mult_Buf[66].Weight_n = Wgt_0_556;
         Mult_Buf[67].Feature_n = FeatureBuf_557;
         Mult_Buf[67].Weight_n = Wgt_0_557;
         Mult_Buf[68].Feature_n = FeatureBuf_558;
         Mult_Buf[68].Weight_n = Wgt_0_558;
         Mult_Buf[69].Feature_n = FeatureBuf_559;
         Mult_Buf[69].Weight_n = Wgt_0_559;
         Mult_Buf[70].Feature_n = FeatureBuf_560;
         Mult_Buf[70].Weight_n = Wgt_0_560;
         Mult_Buf[71].Feature_n = FeatureBuf_561;
         Mult_Buf[71].Weight_n = Wgt_0_561;
         Mult_Buf[72].Feature_n = FeatureBuf_562;
         Mult_Buf[72].Weight_n = Wgt_0_562;
         Mult_Buf[73].Feature_n = FeatureBuf_563;
         Mult_Buf[73].Weight_n = Wgt_0_563;
         Mult_Buf[74].Feature_n = FeatureBuf_564;
         Mult_Buf[74].Weight_n = Wgt_0_564;
         Mult_Buf[75].Feature_n = FeatureBuf_565;
         Mult_Buf[75].Weight_n = Wgt_0_565;
         Mult_Buf[76].Feature_n = FeatureBuf_566;
         Mult_Buf[76].Weight_n = Wgt_0_566;
         Mult_Buf[77].Feature_n = FeatureBuf_567;
         Mult_Buf[77].Weight_n = Wgt_0_567;
         Mult_Buf[78].Feature_n = FeatureBuf_568;
         Mult_Buf[78].Weight_n = Wgt_0_568;
         Mult_Buf[79].Feature_n = FeatureBuf_569;
         Mult_Buf[79].Weight_n = Wgt_0_569;
         Mult_Buf[80].Feature_n = FeatureBuf_570;
         Mult_Buf[80].Weight_n = Wgt_0_570;
         Mult_Buf[81].Feature_n = FeatureBuf_571;
         Mult_Buf[81].Weight_n = Wgt_0_571;
         Mult_Buf[82].Feature_n = FeatureBuf_572;
         Mult_Buf[82].Weight_n = Wgt_0_572;
         Mult_Buf[83].Feature_n = FeatureBuf_573;
         Mult_Buf[83].Weight_n = Wgt_0_573;
         Mult_Buf[84].Feature_n = FeatureBuf_574;
         Mult_Buf[84].Weight_n = Wgt_0_574;
         Mult_Buf[85].Feature_n = FeatureBuf_575;
         Mult_Buf[85].Weight_n = Wgt_0_575;
         Mult_Buf[86].Feature_n = FeatureBuf_576;
         Mult_Buf[86].Weight_n = Wgt_0_576;
         Mult_Buf[87].Feature_n = FeatureBuf_577;
         Mult_Buf[87].Weight_n = Wgt_0_577;
         Mult_Buf[88].Feature_n = FeatureBuf_578;
         Mult_Buf[88].Weight_n = Wgt_0_578;
         Mult_Buf[89].Feature_n = FeatureBuf_579;
         Mult_Buf[89].Weight_n = Wgt_0_579;
         Mult_Buf[90].Feature_n = FeatureBuf_580;
         Mult_Buf[90].Weight_n = Wgt_0_580;
         Mult_Buf[91].Feature_n = FeatureBuf_581;
         Mult_Buf[91].Weight_n = Wgt_0_581;
         Mult_Buf[92].Feature_n = FeatureBuf_582;
         Mult_Buf[92].Weight_n = Wgt_0_582;
         Mult_Buf[93].Feature_n = FeatureBuf_583;
         Mult_Buf[93].Weight_n = Wgt_0_583;
         Mult_Buf[94].Feature_n = FeatureBuf_584;
         Mult_Buf[94].Weight_n = Wgt_0_584;
         Mult_Buf[95].Feature_n = FeatureBuf_585;
         Mult_Buf[95].Weight_n = Wgt_0_585;
         Mult_Buf[96].Feature_n = FeatureBuf_586;
         Mult_Buf[96].Weight_n = Wgt_0_586;
         Mult_Buf[97].Feature_n = FeatureBuf_587;
         Mult_Buf[97].Weight_n = Wgt_0_587;
     end
    8:begin
     nxt_state = 9;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_588;
         Mult_Buf[0].Weight_n = Wgt_0_588;
         Mult_Buf[1].Feature_n = FeatureBuf_589;
         Mult_Buf[1].Weight_n = Wgt_0_589;
         Mult_Buf[2].Feature_n = FeatureBuf_590;
         Mult_Buf[2].Weight_n = Wgt_0_590;
         Mult_Buf[3].Feature_n = FeatureBuf_591;
         Mult_Buf[3].Weight_n = Wgt_0_591;
         Mult_Buf[4].Feature_n = FeatureBuf_592;
         Mult_Buf[4].Weight_n = Wgt_0_592;
         Mult_Buf[5].Feature_n = FeatureBuf_593;
         Mult_Buf[5].Weight_n = Wgt_0_593;
         Mult_Buf[6].Feature_n = FeatureBuf_594;
         Mult_Buf[6].Weight_n = Wgt_0_594;
         Mult_Buf[7].Feature_n = FeatureBuf_595;
         Mult_Buf[7].Weight_n = Wgt_0_595;
         Mult_Buf[8].Feature_n = FeatureBuf_596;
         Mult_Buf[8].Weight_n = Wgt_0_596;
         Mult_Buf[9].Feature_n = FeatureBuf_597;
         Mult_Buf[9].Weight_n = Wgt_0_597;
         Mult_Buf[10].Feature_n = FeatureBuf_598;
         Mult_Buf[10].Weight_n = Wgt_0_598;
         Mult_Buf[11].Feature_n = FeatureBuf_599;
         Mult_Buf[11].Weight_n = Wgt_0_599;
         Mult_Buf[12].Feature_n = FeatureBuf_600;
         Mult_Buf[12].Weight_n = Wgt_0_600;
         Mult_Buf[13].Feature_n = FeatureBuf_601;
         Mult_Buf[13].Weight_n = Wgt_0_601;
         Mult_Buf[14].Feature_n = FeatureBuf_602;
         Mult_Buf[14].Weight_n = Wgt_0_602;
         Mult_Buf[15].Feature_n = FeatureBuf_603;
         Mult_Buf[15].Weight_n = Wgt_0_603;
         Mult_Buf[16].Feature_n = FeatureBuf_604;
         Mult_Buf[16].Weight_n = Wgt_0_604;
         Mult_Buf[17].Feature_n = FeatureBuf_605;
         Mult_Buf[17].Weight_n = Wgt_0_605;
         Mult_Buf[18].Feature_n = FeatureBuf_606;
         Mult_Buf[18].Weight_n = Wgt_0_606;
         Mult_Buf[19].Feature_n = FeatureBuf_607;
         Mult_Buf[19].Weight_n = Wgt_0_607;
         Mult_Buf[20].Feature_n = FeatureBuf_608;
         Mult_Buf[20].Weight_n = Wgt_0_608;
         Mult_Buf[21].Feature_n = FeatureBuf_609;
         Mult_Buf[21].Weight_n = Wgt_0_609;
         Mult_Buf[22].Feature_n = FeatureBuf_610;
         Mult_Buf[22].Weight_n = Wgt_0_610;
         Mult_Buf[23].Feature_n = FeatureBuf_611;
         Mult_Buf[23].Weight_n = Wgt_0_611;
         Mult_Buf[24].Feature_n = FeatureBuf_612;
         Mult_Buf[24].Weight_n = Wgt_0_612;
         Mult_Buf[25].Feature_n = FeatureBuf_613;
         Mult_Buf[25].Weight_n = Wgt_0_613;
         Mult_Buf[26].Feature_n = FeatureBuf_614;
         Mult_Buf[26].Weight_n = Wgt_0_614;
         Mult_Buf[27].Feature_n = FeatureBuf_615;
         Mult_Buf[27].Weight_n = Wgt_0_615;
         Mult_Buf[28].Feature_n = FeatureBuf_616;
         Mult_Buf[28].Weight_n = Wgt_0_616;
         Mult_Buf[29].Feature_n = FeatureBuf_617;
         Mult_Buf[29].Weight_n = Wgt_0_617;
         Mult_Buf[30].Feature_n = FeatureBuf_618;
         Mult_Buf[30].Weight_n = Wgt_0_618;
         Mult_Buf[31].Feature_n = FeatureBuf_619;
         Mult_Buf[31].Weight_n = Wgt_0_619;
         Mult_Buf[32].Feature_n = FeatureBuf_620;
         Mult_Buf[32].Weight_n = Wgt_0_620;
         Mult_Buf[33].Feature_n = FeatureBuf_621;
         Mult_Buf[33].Weight_n = Wgt_0_621;
         Mult_Buf[34].Feature_n = FeatureBuf_622;
         Mult_Buf[34].Weight_n = Wgt_0_622;
         Mult_Buf[35].Feature_n = FeatureBuf_623;
         Mult_Buf[35].Weight_n = Wgt_0_623;
         Mult_Buf[36].Feature_n = FeatureBuf_624;
         Mult_Buf[36].Weight_n = Wgt_0_624;
         Mult_Buf[37].Feature_n = FeatureBuf_625;
         Mult_Buf[37].Weight_n = Wgt_0_625;
         Mult_Buf[38].Feature_n = FeatureBuf_626;
         Mult_Buf[38].Weight_n = Wgt_0_626;
         Mult_Buf[39].Feature_n = FeatureBuf_627;
         Mult_Buf[39].Weight_n = Wgt_0_627;
         Mult_Buf[40].Feature_n = FeatureBuf_628;
         Mult_Buf[40].Weight_n = Wgt_0_628;
         Mult_Buf[41].Feature_n = FeatureBuf_629;
         Mult_Buf[41].Weight_n = Wgt_0_629;
         Mult_Buf[42].Feature_n = FeatureBuf_630;
         Mult_Buf[42].Weight_n = Wgt_0_630;
         Mult_Buf[43].Feature_n = FeatureBuf_631;
         Mult_Buf[43].Weight_n = Wgt_0_631;
         Mult_Buf[44].Feature_n = FeatureBuf_632;
         Mult_Buf[44].Weight_n = Wgt_0_632;
         Mult_Buf[45].Feature_n = FeatureBuf_633;
         Mult_Buf[45].Weight_n = Wgt_0_633;
         Mult_Buf[46].Feature_n = FeatureBuf_634;
         Mult_Buf[46].Weight_n = Wgt_0_634;
         Mult_Buf[47].Feature_n = FeatureBuf_635;
         Mult_Buf[47].Weight_n = Wgt_0_635;
         Mult_Buf[48].Feature_n = FeatureBuf_636;
         Mult_Buf[48].Weight_n = Wgt_0_636;
         Mult_Buf[49].Feature_n = FeatureBuf_637;
         Mult_Buf[49].Weight_n = Wgt_0_637;
         Mult_Buf[50].Feature_n = FeatureBuf_638;
         Mult_Buf[50].Weight_n = Wgt_0_638;
         Mult_Buf[51].Feature_n = FeatureBuf_639;
         Mult_Buf[51].Weight_n = Wgt_0_639;
         Mult_Buf[52].Feature_n = FeatureBuf_640;
         Mult_Buf[52].Weight_n = Wgt_0_640;
         Mult_Buf[53].Feature_n = FeatureBuf_641;
         Mult_Buf[53].Weight_n = Wgt_0_641;
         Mult_Buf[54].Feature_n = FeatureBuf_642;
         Mult_Buf[54].Weight_n = Wgt_0_642;
         Mult_Buf[55].Feature_n = FeatureBuf_643;
         Mult_Buf[55].Weight_n = Wgt_0_643;
         Mult_Buf[56].Feature_n = FeatureBuf_644;
         Mult_Buf[56].Weight_n = Wgt_0_644;
         Mult_Buf[57].Feature_n = FeatureBuf_645;
         Mult_Buf[57].Weight_n = Wgt_0_645;
         Mult_Buf[58].Feature_n = FeatureBuf_646;
         Mult_Buf[58].Weight_n = Wgt_0_646;
         Mult_Buf[59].Feature_n = FeatureBuf_647;
         Mult_Buf[59].Weight_n = Wgt_0_647;
         Mult_Buf[60].Feature_n = FeatureBuf_648;
         Mult_Buf[60].Weight_n = Wgt_0_648;
         Mult_Buf[61].Feature_n = FeatureBuf_649;
         Mult_Buf[61].Weight_n = Wgt_0_649;
         Mult_Buf[62].Feature_n = FeatureBuf_650;
         Mult_Buf[62].Weight_n = Wgt_0_650;
         Mult_Buf[63].Feature_n = FeatureBuf_651;
         Mult_Buf[63].Weight_n = Wgt_0_651;
         Mult_Buf[64].Feature_n = FeatureBuf_652;
         Mult_Buf[64].Weight_n = Wgt_0_652;
         Mult_Buf[65].Feature_n = FeatureBuf_653;
         Mult_Buf[65].Weight_n = Wgt_0_653;
         Mult_Buf[66].Feature_n = FeatureBuf_654;
         Mult_Buf[66].Weight_n = Wgt_0_654;
         Mult_Buf[67].Feature_n = FeatureBuf_655;
         Mult_Buf[67].Weight_n = Wgt_0_655;
         Mult_Buf[68].Feature_n = FeatureBuf_656;
         Mult_Buf[68].Weight_n = Wgt_0_656;
         Mult_Buf[69].Feature_n = FeatureBuf_657;
         Mult_Buf[69].Weight_n = Wgt_0_657;
         Mult_Buf[70].Feature_n = FeatureBuf_658;
         Mult_Buf[70].Weight_n = Wgt_0_658;
         Mult_Buf[71].Feature_n = FeatureBuf_659;
         Mult_Buf[71].Weight_n = Wgt_0_659;
         Mult_Buf[72].Feature_n = FeatureBuf_660;
         Mult_Buf[72].Weight_n = Wgt_0_660;
         Mult_Buf[73].Feature_n = FeatureBuf_661;
         Mult_Buf[73].Weight_n = Wgt_0_661;
         Mult_Buf[74].Feature_n = FeatureBuf_662;
         Mult_Buf[74].Weight_n = Wgt_0_662;
         Mult_Buf[75].Feature_n = FeatureBuf_663;
         Mult_Buf[75].Weight_n = Wgt_0_663;
         Mult_Buf[76].Feature_n = FeatureBuf_664;
         Mult_Buf[76].Weight_n = Wgt_0_664;
         Mult_Buf[77].Feature_n = FeatureBuf_665;
         Mult_Buf[77].Weight_n = Wgt_0_665;
         Mult_Buf[78].Feature_n = FeatureBuf_666;
         Mult_Buf[78].Weight_n = Wgt_0_666;
         Mult_Buf[79].Feature_n = FeatureBuf_667;
         Mult_Buf[79].Weight_n = Wgt_0_667;
         Mult_Buf[80].Feature_n = FeatureBuf_668;
         Mult_Buf[80].Weight_n = Wgt_0_668;
         Mult_Buf[81].Feature_n = FeatureBuf_669;
         Mult_Buf[81].Weight_n = Wgt_0_669;
         Mult_Buf[82].Feature_n = FeatureBuf_670;
         Mult_Buf[82].Weight_n = Wgt_0_670;
         Mult_Buf[83].Feature_n = FeatureBuf_671;
         Mult_Buf[83].Weight_n = Wgt_0_671;
         Mult_Buf[84].Feature_n = FeatureBuf_672;
         Mult_Buf[84].Weight_n = Wgt_0_672;
         Mult_Buf[85].Feature_n = FeatureBuf_673;
         Mult_Buf[85].Weight_n = Wgt_0_673;
         Mult_Buf[86].Feature_n = FeatureBuf_674;
         Mult_Buf[86].Weight_n = Wgt_0_674;
         Mult_Buf[87].Feature_n = FeatureBuf_675;
         Mult_Buf[87].Weight_n = Wgt_0_675;
         Mult_Buf[88].Feature_n = FeatureBuf_676;
         Mult_Buf[88].Weight_n = Wgt_0_676;
         Mult_Buf[89].Feature_n = FeatureBuf_677;
         Mult_Buf[89].Weight_n = Wgt_0_677;
         Mult_Buf[90].Feature_n = FeatureBuf_678;
         Mult_Buf[90].Weight_n = Wgt_0_678;
         Mult_Buf[91].Feature_n = FeatureBuf_679;
         Mult_Buf[91].Weight_n = Wgt_0_679;
         Mult_Buf[92].Feature_n = FeatureBuf_680;
         Mult_Buf[92].Weight_n = Wgt_0_680;
         Mult_Buf[93].Feature_n = FeatureBuf_681;
         Mult_Buf[93].Weight_n = Wgt_0_681;
         Mult_Buf[94].Feature_n = FeatureBuf_682;
         Mult_Buf[94].Weight_n = Wgt_0_682;
         Mult_Buf[95].Feature_n = FeatureBuf_683;
         Mult_Buf[95].Weight_n = Wgt_0_683;
         Mult_Buf[96].Feature_n = FeatureBuf_684;
         Mult_Buf[96].Weight_n = Wgt_0_684;
         Mult_Buf[97].Feature_n = FeatureBuf_685;
         Mult_Buf[97].Weight_n = Wgt_0_685;
     end
    9:begin
     nxt_state = 10;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_686;
         Mult_Buf[0].Weight_n = Wgt_0_686;
         Mult_Buf[1].Feature_n = FeatureBuf_687;
         Mult_Buf[1].Weight_n = Wgt_0_687;
         Mult_Buf[2].Feature_n = FeatureBuf_688;
         Mult_Buf[2].Weight_n = Wgt_0_688;
         Mult_Buf[3].Feature_n = FeatureBuf_689;
         Mult_Buf[3].Weight_n = Wgt_0_689;
         Mult_Buf[4].Feature_n = FeatureBuf_690;
         Mult_Buf[4].Weight_n = Wgt_0_690;
         Mult_Buf[5].Feature_n = FeatureBuf_691;
         Mult_Buf[5].Weight_n = Wgt_0_691;
         Mult_Buf[6].Feature_n = FeatureBuf_692;
         Mult_Buf[6].Weight_n = Wgt_0_692;
         Mult_Buf[7].Feature_n = FeatureBuf_693;
         Mult_Buf[7].Weight_n = Wgt_0_693;
         Mult_Buf[8].Feature_n = FeatureBuf_694;
         Mult_Buf[8].Weight_n = Wgt_0_694;
         Mult_Buf[9].Feature_n = FeatureBuf_695;
         Mult_Buf[9].Weight_n = Wgt_0_695;
         Mult_Buf[10].Feature_n = FeatureBuf_696;
         Mult_Buf[10].Weight_n = Wgt_0_696;
         Mult_Buf[11].Feature_n = FeatureBuf_697;
         Mult_Buf[11].Weight_n = Wgt_0_697;
         Mult_Buf[12].Feature_n = FeatureBuf_698;
         Mult_Buf[12].Weight_n = Wgt_0_698;
         Mult_Buf[13].Feature_n = FeatureBuf_699;
         Mult_Buf[13].Weight_n = Wgt_0_699;
         Mult_Buf[14].Feature_n = FeatureBuf_700;
         Mult_Buf[14].Weight_n = Wgt_0_700;
         Mult_Buf[15].Feature_n = FeatureBuf_701;
         Mult_Buf[15].Weight_n = Wgt_0_701;
         Mult_Buf[16].Feature_n = FeatureBuf_702;
         Mult_Buf[16].Weight_n = Wgt_0_702;
         Mult_Buf[17].Feature_n = FeatureBuf_703;
         Mult_Buf[17].Weight_n = Wgt_0_703;
         Mult_Buf[18].Feature_n = FeatureBuf_704;
         Mult_Buf[18].Weight_n = Wgt_0_704;
         Mult_Buf[19].Feature_n = FeatureBuf_705;
         Mult_Buf[19].Weight_n = Wgt_0_705;
         Mult_Buf[20].Feature_n = FeatureBuf_706;
         Mult_Buf[20].Weight_n = Wgt_0_706;
         Mult_Buf[21].Feature_n = FeatureBuf_707;
         Mult_Buf[21].Weight_n = Wgt_0_707;
         Mult_Buf[22].Feature_n = FeatureBuf_708;
         Mult_Buf[22].Weight_n = Wgt_0_708;
         Mult_Buf[23].Feature_n = FeatureBuf_709;
         Mult_Buf[23].Weight_n = Wgt_0_709;
         Mult_Buf[24].Feature_n = FeatureBuf_710;
         Mult_Buf[24].Weight_n = Wgt_0_710;
         Mult_Buf[25].Feature_n = FeatureBuf_711;
         Mult_Buf[25].Weight_n = Wgt_0_711;
         Mult_Buf[26].Feature_n = FeatureBuf_712;
         Mult_Buf[26].Weight_n = Wgt_0_712;
         Mult_Buf[27].Feature_n = FeatureBuf_713;
         Mult_Buf[27].Weight_n = Wgt_0_713;
         Mult_Buf[28].Feature_n = FeatureBuf_714;
         Mult_Buf[28].Weight_n = Wgt_0_714;
         Mult_Buf[29].Feature_n = FeatureBuf_715;
         Mult_Buf[29].Weight_n = Wgt_0_715;
         Mult_Buf[30].Feature_n = FeatureBuf_716;
         Mult_Buf[30].Weight_n = Wgt_0_716;
         Mult_Buf[31].Feature_n = FeatureBuf_717;
         Mult_Buf[31].Weight_n = Wgt_0_717;
         Mult_Buf[32].Feature_n = FeatureBuf_718;
         Mult_Buf[32].Weight_n = Wgt_0_718;
         Mult_Buf[33].Feature_n = FeatureBuf_719;
         Mult_Buf[33].Weight_n = Wgt_0_719;
         Mult_Buf[34].Feature_n = FeatureBuf_720;
         Mult_Buf[34].Weight_n = Wgt_0_720;
         Mult_Buf[35].Feature_n = FeatureBuf_721;
         Mult_Buf[35].Weight_n = Wgt_0_721;
         Mult_Buf[36].Feature_n = FeatureBuf_722;
         Mult_Buf[36].Weight_n = Wgt_0_722;
         Mult_Buf[37].Feature_n = FeatureBuf_723;
         Mult_Buf[37].Weight_n = Wgt_0_723;
         Mult_Buf[38].Feature_n = FeatureBuf_724;
         Mult_Buf[38].Weight_n = Wgt_0_724;
         Mult_Buf[39].Feature_n = FeatureBuf_725;
         Mult_Buf[39].Weight_n = Wgt_0_725;
         Mult_Buf[40].Feature_n = FeatureBuf_726;
         Mult_Buf[40].Weight_n = Wgt_0_726;
         Mult_Buf[41].Feature_n = FeatureBuf_727;
         Mult_Buf[41].Weight_n = Wgt_0_727;
         Mult_Buf[42].Feature_n = FeatureBuf_728;
         Mult_Buf[42].Weight_n = Wgt_0_728;
         Mult_Buf[43].Feature_n = FeatureBuf_729;
         Mult_Buf[43].Weight_n = Wgt_0_729;
         Mult_Buf[44].Feature_n = FeatureBuf_730;
         Mult_Buf[44].Weight_n = Wgt_0_730;
         Mult_Buf[45].Feature_n = FeatureBuf_731;
         Mult_Buf[45].Weight_n = Wgt_0_731;
         Mult_Buf[46].Feature_n = FeatureBuf_732;
         Mult_Buf[46].Weight_n = Wgt_0_732;
         Mult_Buf[47].Feature_n = FeatureBuf_733;
         Mult_Buf[47].Weight_n = Wgt_0_733;
         Mult_Buf[48].Feature_n = FeatureBuf_734;
         Mult_Buf[48].Weight_n = Wgt_0_734;
         Mult_Buf[49].Feature_n = FeatureBuf_735;
         Mult_Buf[49].Weight_n = Wgt_0_735;
         Mult_Buf[50].Feature_n = FeatureBuf_736;
         Mult_Buf[50].Weight_n = Wgt_0_736;
         Mult_Buf[51].Feature_n = FeatureBuf_737;
         Mult_Buf[51].Weight_n = Wgt_0_737;
         Mult_Buf[52].Feature_n = FeatureBuf_738;
         Mult_Buf[52].Weight_n = Wgt_0_738;
         Mult_Buf[53].Feature_n = FeatureBuf_739;
         Mult_Buf[53].Weight_n = Wgt_0_739;
         Mult_Buf[54].Feature_n = FeatureBuf_740;
         Mult_Buf[54].Weight_n = Wgt_0_740;
         Mult_Buf[55].Feature_n = FeatureBuf_741;
         Mult_Buf[55].Weight_n = Wgt_0_741;
         Mult_Buf[56].Feature_n = FeatureBuf_742;
         Mult_Buf[56].Weight_n = Wgt_0_742;
         Mult_Buf[57].Feature_n = FeatureBuf_743;
         Mult_Buf[57].Weight_n = Wgt_0_743;
         Mult_Buf[58].Feature_n = FeatureBuf_744;
         Mult_Buf[58].Weight_n = Wgt_0_744;
         Mult_Buf[59].Feature_n = FeatureBuf_745;
         Mult_Buf[59].Weight_n = Wgt_0_745;
         Mult_Buf[60].Feature_n = FeatureBuf_746;
         Mult_Buf[60].Weight_n = Wgt_0_746;
         Mult_Buf[61].Feature_n = FeatureBuf_747;
         Mult_Buf[61].Weight_n = Wgt_0_747;
         Mult_Buf[62].Feature_n = FeatureBuf_748;
         Mult_Buf[62].Weight_n = Wgt_0_748;
         Mult_Buf[63].Feature_n = FeatureBuf_749;
         Mult_Buf[63].Weight_n = Wgt_0_749;
         Mult_Buf[64].Feature_n = FeatureBuf_750;
         Mult_Buf[64].Weight_n = Wgt_0_750;
         Mult_Buf[65].Feature_n = FeatureBuf_751;
         Mult_Buf[65].Weight_n = Wgt_0_751;
         Mult_Buf[66].Feature_n = FeatureBuf_752;
         Mult_Buf[66].Weight_n = Wgt_0_752;
         Mult_Buf[67].Feature_n = FeatureBuf_753;
         Mult_Buf[67].Weight_n = Wgt_0_753;
         Mult_Buf[68].Feature_n = FeatureBuf_754;
         Mult_Buf[68].Weight_n = Wgt_0_754;
         Mult_Buf[69].Feature_n = FeatureBuf_755;
         Mult_Buf[69].Weight_n = Wgt_0_755;
         Mult_Buf[70].Feature_n = FeatureBuf_756;
         Mult_Buf[70].Weight_n = Wgt_0_756;
         Mult_Buf[71].Feature_n = FeatureBuf_757;
         Mult_Buf[71].Weight_n = Wgt_0_757;
         Mult_Buf[72].Feature_n = FeatureBuf_758;
         Mult_Buf[72].Weight_n = Wgt_0_758;
         Mult_Buf[73].Feature_n = FeatureBuf_759;
         Mult_Buf[73].Weight_n = Wgt_0_759;
         Mult_Buf[74].Feature_n = FeatureBuf_760;
         Mult_Buf[74].Weight_n = Wgt_0_760;
         Mult_Buf[75].Feature_n = FeatureBuf_761;
         Mult_Buf[75].Weight_n = Wgt_0_761;
         Mult_Buf[76].Feature_n = FeatureBuf_762;
         Mult_Buf[76].Weight_n = Wgt_0_762;
         Mult_Buf[77].Feature_n = FeatureBuf_763;
         Mult_Buf[77].Weight_n = Wgt_0_763;
         Mult_Buf[78].Feature_n = FeatureBuf_764;
         Mult_Buf[78].Weight_n = Wgt_0_764;
         Mult_Buf[79].Feature_n = FeatureBuf_765;
         Mult_Buf[79].Weight_n = Wgt_0_765;
         Mult_Buf[80].Feature_n = FeatureBuf_766;
         Mult_Buf[80].Weight_n = Wgt_0_766;
         Mult_Buf[81].Feature_n = FeatureBuf_767;
         Mult_Buf[81].Weight_n = Wgt_0_767;
         Mult_Buf[82].Feature_n = FeatureBuf_768;
         Mult_Buf[82].Weight_n = Wgt_0_768;
         Mult_Buf[83].Feature_n = FeatureBuf_769;
         Mult_Buf[83].Weight_n = Wgt_0_769;
         Mult_Buf[84].Feature_n = FeatureBuf_770;
         Mult_Buf[84].Weight_n = Wgt_0_770;
         Mult_Buf[85].Feature_n = FeatureBuf_771;
         Mult_Buf[85].Weight_n = Wgt_0_771;
         Mult_Buf[86].Feature_n = FeatureBuf_772;
         Mult_Buf[86].Weight_n = Wgt_0_772;
         Mult_Buf[87].Feature_n = FeatureBuf_773;
         Mult_Buf[87].Weight_n = Wgt_0_773;
         Mult_Buf[88].Feature_n = FeatureBuf_774;
         Mult_Buf[88].Weight_n = Wgt_0_774;
         Mult_Buf[89].Feature_n = FeatureBuf_775;
         Mult_Buf[89].Weight_n = Wgt_0_775;
         Mult_Buf[90].Feature_n = FeatureBuf_776;
         Mult_Buf[90].Weight_n = Wgt_0_776;
         Mult_Buf[91].Feature_n = FeatureBuf_777;
         Mult_Buf[91].Weight_n = Wgt_0_777;
         Mult_Buf[92].Feature_n = FeatureBuf_778;
         Mult_Buf[92].Weight_n = Wgt_0_778;
         Mult_Buf[93].Feature_n = FeatureBuf_779;
         Mult_Buf[93].Weight_n = Wgt_0_779;
         Mult_Buf[94].Feature_n = FeatureBuf_780;
         Mult_Buf[94].Weight_n = Wgt_0_780;
         Mult_Buf[95].Feature_n = FeatureBuf_781;
         Mult_Buf[95].Weight_n = Wgt_0_781;
         Mult_Buf[96].Feature_n = FeatureBuf_782;
         Mult_Buf[96].Weight_n = Wgt_0_782;
         Mult_Buf[97].Feature_n = FeatureBuf_783;
         Mult_Buf[97].Weight_n = Wgt_0_783;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     end
    10:begin
     nxt_state = 11;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_0;
         Mult_Buf[0].Weight_n = Wgt_1_0;
         Mult_Buf[1].Feature_n = FeatureBuf_1;
         Mult_Buf[1].Weight_n = Wgt_1_1;
         Mult_Buf[2].Feature_n = FeatureBuf_2;
         Mult_Buf[2].Weight_n = Wgt_1_2;
         Mult_Buf[3].Feature_n = FeatureBuf_3;
         Mult_Buf[3].Weight_n = Wgt_1_3;
         Mult_Buf[4].Feature_n = FeatureBuf_4;
         Mult_Buf[4].Weight_n = Wgt_1_4;
         Mult_Buf[5].Feature_n = FeatureBuf_5;
         Mult_Buf[5].Weight_n = Wgt_1_5;
         Mult_Buf[6].Feature_n = FeatureBuf_6;
         Mult_Buf[6].Weight_n = Wgt_1_6;
         Mult_Buf[7].Feature_n = FeatureBuf_7;
         Mult_Buf[7].Weight_n = Wgt_1_7;
         Mult_Buf[8].Feature_n = FeatureBuf_8;
         Mult_Buf[8].Weight_n = Wgt_1_8;
         Mult_Buf[9].Feature_n = FeatureBuf_9;
         Mult_Buf[9].Weight_n = Wgt_1_9;
         Mult_Buf[10].Feature_n = FeatureBuf_10;
         Mult_Buf[10].Weight_n = Wgt_1_10;
         Mult_Buf[11].Feature_n = FeatureBuf_11;
         Mult_Buf[11].Weight_n = Wgt_1_11;
         Mult_Buf[12].Feature_n = FeatureBuf_12;
         Mult_Buf[12].Weight_n = Wgt_1_12;
         Mult_Buf[13].Feature_n = FeatureBuf_13;
         Mult_Buf[13].Weight_n = Wgt_1_13;
         Mult_Buf[14].Feature_n = FeatureBuf_14;
         Mult_Buf[14].Weight_n = Wgt_1_14;
         Mult_Buf[15].Feature_n = FeatureBuf_15;
         Mult_Buf[15].Weight_n = Wgt_1_15;
         Mult_Buf[16].Feature_n = FeatureBuf_16;
         Mult_Buf[16].Weight_n = Wgt_1_16;
         Mult_Buf[17].Feature_n = FeatureBuf_17;
         Mult_Buf[17].Weight_n = Wgt_1_17;
         Mult_Buf[18].Feature_n = FeatureBuf_18;
         Mult_Buf[18].Weight_n = Wgt_1_18;
         Mult_Buf[19].Feature_n = FeatureBuf_19;
         Mult_Buf[19].Weight_n = Wgt_1_19;
         Mult_Buf[20].Feature_n = FeatureBuf_20;
         Mult_Buf[20].Weight_n = Wgt_1_20;
         Mult_Buf[21].Feature_n = FeatureBuf_21;
         Mult_Buf[21].Weight_n = Wgt_1_21;
         Mult_Buf[22].Feature_n = FeatureBuf_22;
         Mult_Buf[22].Weight_n = Wgt_1_22;
         Mult_Buf[23].Feature_n = FeatureBuf_23;
         Mult_Buf[23].Weight_n = Wgt_1_23;
         Mult_Buf[24].Feature_n = FeatureBuf_24;
         Mult_Buf[24].Weight_n = Wgt_1_24;
         Mult_Buf[25].Feature_n = FeatureBuf_25;
         Mult_Buf[25].Weight_n = Wgt_1_25;
         Mult_Buf[26].Feature_n = FeatureBuf_26;
         Mult_Buf[26].Weight_n = Wgt_1_26;
         Mult_Buf[27].Feature_n = FeatureBuf_27;
         Mult_Buf[27].Weight_n = Wgt_1_27;
         Mult_Buf[28].Feature_n = FeatureBuf_28;
         Mult_Buf[28].Weight_n = Wgt_1_28;
         Mult_Buf[29].Feature_n = FeatureBuf_29;
         Mult_Buf[29].Weight_n = Wgt_1_29;
         Mult_Buf[30].Feature_n = FeatureBuf_30;
         Mult_Buf[30].Weight_n = Wgt_1_30;
         Mult_Buf[31].Feature_n = FeatureBuf_31;
         Mult_Buf[31].Weight_n = Wgt_1_31;
         Mult_Buf[32].Feature_n = FeatureBuf_32;
         Mult_Buf[32].Weight_n = Wgt_1_32;
         Mult_Buf[33].Feature_n = FeatureBuf_33;
         Mult_Buf[33].Weight_n = Wgt_1_33;
         Mult_Buf[34].Feature_n = FeatureBuf_34;
         Mult_Buf[34].Weight_n = Wgt_1_34;
         Mult_Buf[35].Feature_n = FeatureBuf_35;
         Mult_Buf[35].Weight_n = Wgt_1_35;
         Mult_Buf[36].Feature_n = FeatureBuf_36;
         Mult_Buf[36].Weight_n = Wgt_1_36;
         Mult_Buf[37].Feature_n = FeatureBuf_37;
         Mult_Buf[37].Weight_n = Wgt_1_37;
         Mult_Buf[38].Feature_n = FeatureBuf_38;
         Mult_Buf[38].Weight_n = Wgt_1_38;
         Mult_Buf[39].Feature_n = FeatureBuf_39;
         Mult_Buf[39].Weight_n = Wgt_1_39;
         Mult_Buf[40].Feature_n = FeatureBuf_40;
         Mult_Buf[40].Weight_n = Wgt_1_40;
         Mult_Buf[41].Feature_n = FeatureBuf_41;
         Mult_Buf[41].Weight_n = Wgt_1_41;
         Mult_Buf[42].Feature_n = FeatureBuf_42;
         Mult_Buf[42].Weight_n = Wgt_1_42;
         Mult_Buf[43].Feature_n = FeatureBuf_43;
         Mult_Buf[43].Weight_n = Wgt_1_43;
         Mult_Buf[44].Feature_n = FeatureBuf_44;
         Mult_Buf[44].Weight_n = Wgt_1_44;
         Mult_Buf[45].Feature_n = FeatureBuf_45;
         Mult_Buf[45].Weight_n = Wgt_1_45;
         Mult_Buf[46].Feature_n = FeatureBuf_46;
         Mult_Buf[46].Weight_n = Wgt_1_46;
         Mult_Buf[47].Feature_n = FeatureBuf_47;
         Mult_Buf[47].Weight_n = Wgt_1_47;
         Mult_Buf[48].Feature_n = FeatureBuf_48;
         Mult_Buf[48].Weight_n = Wgt_1_48;
         Mult_Buf[49].Feature_n = FeatureBuf_49;
         Mult_Buf[49].Weight_n = Wgt_1_49;
         Mult_Buf[50].Feature_n = FeatureBuf_50;
         Mult_Buf[50].Weight_n = Wgt_1_50;
         Mult_Buf[51].Feature_n = FeatureBuf_51;
         Mult_Buf[51].Weight_n = Wgt_1_51;
         Mult_Buf[52].Feature_n = FeatureBuf_52;
         Mult_Buf[52].Weight_n = Wgt_1_52;
         Mult_Buf[53].Feature_n = FeatureBuf_53;
         Mult_Buf[53].Weight_n = Wgt_1_53;
         Mult_Buf[54].Feature_n = FeatureBuf_54;
         Mult_Buf[54].Weight_n = Wgt_1_54;
         Mult_Buf[55].Feature_n = FeatureBuf_55;
         Mult_Buf[55].Weight_n = Wgt_1_55;
         Mult_Buf[56].Feature_n = FeatureBuf_56;
         Mult_Buf[56].Weight_n = Wgt_1_56;
         Mult_Buf[57].Feature_n = FeatureBuf_57;
         Mult_Buf[57].Weight_n = Wgt_1_57;
         Mult_Buf[58].Feature_n = FeatureBuf_58;
         Mult_Buf[58].Weight_n = Wgt_1_58;
         Mult_Buf[59].Feature_n = FeatureBuf_59;
         Mult_Buf[59].Weight_n = Wgt_1_59;
         Mult_Buf[60].Feature_n = FeatureBuf_60;
         Mult_Buf[60].Weight_n = Wgt_1_60;
         Mult_Buf[61].Feature_n = FeatureBuf_61;
         Mult_Buf[61].Weight_n = Wgt_1_61;
         Mult_Buf[62].Feature_n = FeatureBuf_62;
         Mult_Buf[62].Weight_n = Wgt_1_62;
         Mult_Buf[63].Feature_n = FeatureBuf_63;
         Mult_Buf[63].Weight_n = Wgt_1_63;
         Mult_Buf[64].Feature_n = FeatureBuf_64;
         Mult_Buf[64].Weight_n = Wgt_1_64;
         Mult_Buf[65].Feature_n = FeatureBuf_65;
         Mult_Buf[65].Weight_n = Wgt_1_65;
         Mult_Buf[66].Feature_n = FeatureBuf_66;
         Mult_Buf[66].Weight_n = Wgt_1_66;
         Mult_Buf[67].Feature_n = FeatureBuf_67;
         Mult_Buf[67].Weight_n = Wgt_1_67;
         Mult_Buf[68].Feature_n = FeatureBuf_68;
         Mult_Buf[68].Weight_n = Wgt_1_68;
         Mult_Buf[69].Feature_n = FeatureBuf_69;
         Mult_Buf[69].Weight_n = Wgt_1_69;
         Mult_Buf[70].Feature_n = FeatureBuf_70;
         Mult_Buf[70].Weight_n = Wgt_1_70;
         Mult_Buf[71].Feature_n = FeatureBuf_71;
         Mult_Buf[71].Weight_n = Wgt_1_71;
         Mult_Buf[72].Feature_n = FeatureBuf_72;
         Mult_Buf[72].Weight_n = Wgt_1_72;
         Mult_Buf[73].Feature_n = FeatureBuf_73;
         Mult_Buf[73].Weight_n = Wgt_1_73;
         Mult_Buf[74].Feature_n = FeatureBuf_74;
         Mult_Buf[74].Weight_n = Wgt_1_74;
         Mult_Buf[75].Feature_n = FeatureBuf_75;
         Mult_Buf[75].Weight_n = Wgt_1_75;
         Mult_Buf[76].Feature_n = FeatureBuf_76;
         Mult_Buf[76].Weight_n = Wgt_1_76;
         Mult_Buf[77].Feature_n = FeatureBuf_77;
         Mult_Buf[77].Weight_n = Wgt_1_77;
         Mult_Buf[78].Feature_n = FeatureBuf_78;
         Mult_Buf[78].Weight_n = Wgt_1_78;
         Mult_Buf[79].Feature_n = FeatureBuf_79;
         Mult_Buf[79].Weight_n = Wgt_1_79;
         Mult_Buf[80].Feature_n = FeatureBuf_80;
         Mult_Buf[80].Weight_n = Wgt_1_80;
         Mult_Buf[81].Feature_n = FeatureBuf_81;
         Mult_Buf[81].Weight_n = Wgt_1_81;
         Mult_Buf[82].Feature_n = FeatureBuf_82;
         Mult_Buf[82].Weight_n = Wgt_1_82;
         Mult_Buf[83].Feature_n = FeatureBuf_83;
         Mult_Buf[83].Weight_n = Wgt_1_83;
         Mult_Buf[84].Feature_n = FeatureBuf_84;
         Mult_Buf[84].Weight_n = Wgt_1_84;
         Mult_Buf[85].Feature_n = FeatureBuf_85;
         Mult_Buf[85].Weight_n = Wgt_1_85;
         Mult_Buf[86].Feature_n = FeatureBuf_86;
         Mult_Buf[86].Weight_n = Wgt_1_86;
         Mult_Buf[87].Feature_n = FeatureBuf_87;
         Mult_Buf[87].Weight_n = Wgt_1_87;
         Mult_Buf[88].Feature_n = FeatureBuf_88;
         Mult_Buf[88].Weight_n = Wgt_1_88;
         Mult_Buf[89].Feature_n = FeatureBuf_89;
         Mult_Buf[89].Weight_n = Wgt_1_89;
         Mult_Buf[90].Feature_n = FeatureBuf_90;
         Mult_Buf[90].Weight_n = Wgt_1_90;
         Mult_Buf[91].Feature_n = FeatureBuf_91;
         Mult_Buf[91].Weight_n = Wgt_1_91;
         Mult_Buf[92].Feature_n = FeatureBuf_92;
         Mult_Buf[92].Weight_n = Wgt_1_92;
         Mult_Buf[93].Feature_n = FeatureBuf_93;
         Mult_Buf[93].Weight_n = Wgt_1_93;
         Mult_Buf[94].Feature_n = FeatureBuf_94;
         Mult_Buf[94].Weight_n = Wgt_1_94;
         Mult_Buf[95].Feature_n = FeatureBuf_95;
         Mult_Buf[95].Weight_n = Wgt_1_95;
         Mult_Buf[96].Feature_n = FeatureBuf_96;
         Mult_Buf[96].Weight_n = Wgt_1_96;
         Mult_Buf[97].Feature_n = FeatureBuf_97;
         Mult_Buf[97].Weight_n = Wgt_1_97;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     end
    11:begin
     nxt_state = 12;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_98;
         Mult_Buf[0].Weight_n = Wgt_1_98;
         Mult_Buf[1].Feature_n = FeatureBuf_99;
         Mult_Buf[1].Weight_n = Wgt_1_99;
         Mult_Buf[2].Feature_n = FeatureBuf_100;
         Mult_Buf[2].Weight_n = Wgt_1_100;
         Mult_Buf[3].Feature_n = FeatureBuf_101;
         Mult_Buf[3].Weight_n = Wgt_1_101;
         Mult_Buf[4].Feature_n = FeatureBuf_102;
         Mult_Buf[4].Weight_n = Wgt_1_102;
         Mult_Buf[5].Feature_n = FeatureBuf_103;
         Mult_Buf[5].Weight_n = Wgt_1_103;
         Mult_Buf[6].Feature_n = FeatureBuf_104;
         Mult_Buf[6].Weight_n = Wgt_1_104;
         Mult_Buf[7].Feature_n = FeatureBuf_105;
         Mult_Buf[7].Weight_n = Wgt_1_105;
         Mult_Buf[8].Feature_n = FeatureBuf_106;
         Mult_Buf[8].Weight_n = Wgt_1_106;
         Mult_Buf[9].Feature_n = FeatureBuf_107;
         Mult_Buf[9].Weight_n = Wgt_1_107;
         Mult_Buf[10].Feature_n = FeatureBuf_108;
         Mult_Buf[10].Weight_n = Wgt_1_108;
         Mult_Buf[11].Feature_n = FeatureBuf_109;
         Mult_Buf[11].Weight_n = Wgt_1_109;
         Mult_Buf[12].Feature_n = FeatureBuf_110;
         Mult_Buf[12].Weight_n = Wgt_1_110;
         Mult_Buf[13].Feature_n = FeatureBuf_111;
         Mult_Buf[13].Weight_n = Wgt_1_111;
         Mult_Buf[14].Feature_n = FeatureBuf_112;
         Mult_Buf[14].Weight_n = Wgt_1_112;
         Mult_Buf[15].Feature_n = FeatureBuf_113;
         Mult_Buf[15].Weight_n = Wgt_1_113;
         Mult_Buf[16].Feature_n = FeatureBuf_114;
         Mult_Buf[16].Weight_n = Wgt_1_114;
         Mult_Buf[17].Feature_n = FeatureBuf_115;
         Mult_Buf[17].Weight_n = Wgt_1_115;
         Mult_Buf[18].Feature_n = FeatureBuf_116;
         Mult_Buf[18].Weight_n = Wgt_1_116;
         Mult_Buf[19].Feature_n = FeatureBuf_117;
         Mult_Buf[19].Weight_n = Wgt_1_117;
         Mult_Buf[20].Feature_n = FeatureBuf_118;
         Mult_Buf[20].Weight_n = Wgt_1_118;
         Mult_Buf[21].Feature_n = FeatureBuf_119;
         Mult_Buf[21].Weight_n = Wgt_1_119;
         Mult_Buf[22].Feature_n = FeatureBuf_120;
         Mult_Buf[22].Weight_n = Wgt_1_120;
         Mult_Buf[23].Feature_n = FeatureBuf_121;
         Mult_Buf[23].Weight_n = Wgt_1_121;
         Mult_Buf[24].Feature_n = FeatureBuf_122;
         Mult_Buf[24].Weight_n = Wgt_1_122;
         Mult_Buf[25].Feature_n = FeatureBuf_123;
         Mult_Buf[25].Weight_n = Wgt_1_123;
         Mult_Buf[26].Feature_n = FeatureBuf_124;
         Mult_Buf[26].Weight_n = Wgt_1_124;
         Mult_Buf[27].Feature_n = FeatureBuf_125;
         Mult_Buf[27].Weight_n = Wgt_1_125;
         Mult_Buf[28].Feature_n = FeatureBuf_126;
         Mult_Buf[28].Weight_n = Wgt_1_126;
         Mult_Buf[29].Feature_n = FeatureBuf_127;
         Mult_Buf[29].Weight_n = Wgt_1_127;
         Mult_Buf[30].Feature_n = FeatureBuf_128;
         Mult_Buf[30].Weight_n = Wgt_1_128;
         Mult_Buf[31].Feature_n = FeatureBuf_129;
         Mult_Buf[31].Weight_n = Wgt_1_129;
         Mult_Buf[32].Feature_n = FeatureBuf_130;
         Mult_Buf[32].Weight_n = Wgt_1_130;
         Mult_Buf[33].Feature_n = FeatureBuf_131;
         Mult_Buf[33].Weight_n = Wgt_1_131;
         Mult_Buf[34].Feature_n = FeatureBuf_132;
         Mult_Buf[34].Weight_n = Wgt_1_132;
         Mult_Buf[35].Feature_n = FeatureBuf_133;
         Mult_Buf[35].Weight_n = Wgt_1_133;
         Mult_Buf[36].Feature_n = FeatureBuf_134;
         Mult_Buf[36].Weight_n = Wgt_1_134;
         Mult_Buf[37].Feature_n = FeatureBuf_135;
         Mult_Buf[37].Weight_n = Wgt_1_135;
         Mult_Buf[38].Feature_n = FeatureBuf_136;
         Mult_Buf[38].Weight_n = Wgt_1_136;
         Mult_Buf[39].Feature_n = FeatureBuf_137;
         Mult_Buf[39].Weight_n = Wgt_1_137;
         Mult_Buf[40].Feature_n = FeatureBuf_138;
         Mult_Buf[40].Weight_n = Wgt_1_138;
         Mult_Buf[41].Feature_n = FeatureBuf_139;
         Mult_Buf[41].Weight_n = Wgt_1_139;
         Mult_Buf[42].Feature_n = FeatureBuf_140;
         Mult_Buf[42].Weight_n = Wgt_1_140;
         Mult_Buf[43].Feature_n = FeatureBuf_141;
         Mult_Buf[43].Weight_n = Wgt_1_141;
         Mult_Buf[44].Feature_n = FeatureBuf_142;
         Mult_Buf[44].Weight_n = Wgt_1_142;
         Mult_Buf[45].Feature_n = FeatureBuf_143;
         Mult_Buf[45].Weight_n = Wgt_1_143;
         Mult_Buf[46].Feature_n = FeatureBuf_144;
         Mult_Buf[46].Weight_n = Wgt_1_144;
         Mult_Buf[47].Feature_n = FeatureBuf_145;
         Mult_Buf[47].Weight_n = Wgt_1_145;
         Mult_Buf[48].Feature_n = FeatureBuf_146;
         Mult_Buf[48].Weight_n = Wgt_1_146;
         Mult_Buf[49].Feature_n = FeatureBuf_147;
         Mult_Buf[49].Weight_n = Wgt_1_147;
         Mult_Buf[50].Feature_n = FeatureBuf_148;
         Mult_Buf[50].Weight_n = Wgt_1_148;
         Mult_Buf[51].Feature_n = FeatureBuf_149;
         Mult_Buf[51].Weight_n = Wgt_1_149;
         Mult_Buf[52].Feature_n = FeatureBuf_150;
         Mult_Buf[52].Weight_n = Wgt_1_150;
         Mult_Buf[53].Feature_n = FeatureBuf_151;
         Mult_Buf[53].Weight_n = Wgt_1_151;
         Mult_Buf[54].Feature_n = FeatureBuf_152;
         Mult_Buf[54].Weight_n = Wgt_1_152;
         Mult_Buf[55].Feature_n = FeatureBuf_153;
         Mult_Buf[55].Weight_n = Wgt_1_153;
         Mult_Buf[56].Feature_n = FeatureBuf_154;
         Mult_Buf[56].Weight_n = Wgt_1_154;
         Mult_Buf[57].Feature_n = FeatureBuf_155;
         Mult_Buf[57].Weight_n = Wgt_1_155;
         Mult_Buf[58].Feature_n = FeatureBuf_156;
         Mult_Buf[58].Weight_n = Wgt_1_156;
         Mult_Buf[59].Feature_n = FeatureBuf_157;
         Mult_Buf[59].Weight_n = Wgt_1_157;
         Mult_Buf[60].Feature_n = FeatureBuf_158;
         Mult_Buf[60].Weight_n = Wgt_1_158;
         Mult_Buf[61].Feature_n = FeatureBuf_159;
         Mult_Buf[61].Weight_n = Wgt_1_159;
         Mult_Buf[62].Feature_n = FeatureBuf_160;
         Mult_Buf[62].Weight_n = Wgt_1_160;
         Mult_Buf[63].Feature_n = FeatureBuf_161;
         Mult_Buf[63].Weight_n = Wgt_1_161;
         Mult_Buf[64].Feature_n = FeatureBuf_162;
         Mult_Buf[64].Weight_n = Wgt_1_162;
         Mult_Buf[65].Feature_n = FeatureBuf_163;
         Mult_Buf[65].Weight_n = Wgt_1_163;
         Mult_Buf[66].Feature_n = FeatureBuf_164;
         Mult_Buf[66].Weight_n = Wgt_1_164;
         Mult_Buf[67].Feature_n = FeatureBuf_165;
         Mult_Buf[67].Weight_n = Wgt_1_165;
         Mult_Buf[68].Feature_n = FeatureBuf_166;
         Mult_Buf[68].Weight_n = Wgt_1_166;
         Mult_Buf[69].Feature_n = FeatureBuf_167;
         Mult_Buf[69].Weight_n = Wgt_1_167;
         Mult_Buf[70].Feature_n = FeatureBuf_168;
         Mult_Buf[70].Weight_n = Wgt_1_168;
         Mult_Buf[71].Feature_n = FeatureBuf_169;
         Mult_Buf[71].Weight_n = Wgt_1_169;
         Mult_Buf[72].Feature_n = FeatureBuf_170;
         Mult_Buf[72].Weight_n = Wgt_1_170;
         Mult_Buf[73].Feature_n = FeatureBuf_171;
         Mult_Buf[73].Weight_n = Wgt_1_171;
         Mult_Buf[74].Feature_n = FeatureBuf_172;
         Mult_Buf[74].Weight_n = Wgt_1_172;
         Mult_Buf[75].Feature_n = FeatureBuf_173;
         Mult_Buf[75].Weight_n = Wgt_1_173;
         Mult_Buf[76].Feature_n = FeatureBuf_174;
         Mult_Buf[76].Weight_n = Wgt_1_174;
         Mult_Buf[77].Feature_n = FeatureBuf_175;
         Mult_Buf[77].Weight_n = Wgt_1_175;
         Mult_Buf[78].Feature_n = FeatureBuf_176;
         Mult_Buf[78].Weight_n = Wgt_1_176;
         Mult_Buf[79].Feature_n = FeatureBuf_177;
         Mult_Buf[79].Weight_n = Wgt_1_177;
         Mult_Buf[80].Feature_n = FeatureBuf_178;
         Mult_Buf[80].Weight_n = Wgt_1_178;
         Mult_Buf[81].Feature_n = FeatureBuf_179;
         Mult_Buf[81].Weight_n = Wgt_1_179;
         Mult_Buf[82].Feature_n = FeatureBuf_180;
         Mult_Buf[82].Weight_n = Wgt_1_180;
         Mult_Buf[83].Feature_n = FeatureBuf_181;
         Mult_Buf[83].Weight_n = Wgt_1_181;
         Mult_Buf[84].Feature_n = FeatureBuf_182;
         Mult_Buf[84].Weight_n = Wgt_1_182;
         Mult_Buf[85].Feature_n = FeatureBuf_183;
         Mult_Buf[85].Weight_n = Wgt_1_183;
         Mult_Buf[86].Feature_n = FeatureBuf_184;
         Mult_Buf[86].Weight_n = Wgt_1_184;
         Mult_Buf[87].Feature_n = FeatureBuf_185;
         Mult_Buf[87].Weight_n = Wgt_1_185;
         Mult_Buf[88].Feature_n = FeatureBuf_186;
         Mult_Buf[88].Weight_n = Wgt_1_186;
         Mult_Buf[89].Feature_n = FeatureBuf_187;
         Mult_Buf[89].Weight_n = Wgt_1_187;
         Mult_Buf[90].Feature_n = FeatureBuf_188;
         Mult_Buf[90].Weight_n = Wgt_1_188;
         Mult_Buf[91].Feature_n = FeatureBuf_189;
         Mult_Buf[91].Weight_n = Wgt_1_189;
         Mult_Buf[92].Feature_n = FeatureBuf_190;
         Mult_Buf[92].Weight_n = Wgt_1_190;
         Mult_Buf[93].Feature_n = FeatureBuf_191;
         Mult_Buf[93].Weight_n = Wgt_1_191;
         Mult_Buf[94].Feature_n = FeatureBuf_192;
         Mult_Buf[94].Weight_n = Wgt_1_192;
         Mult_Buf[95].Feature_n = FeatureBuf_193;
         Mult_Buf[95].Weight_n = Wgt_1_193;
         Mult_Buf[96].Feature_n = FeatureBuf_194;
         Mult_Buf[96].Weight_n = Wgt_1_194;
         Mult_Buf[97].Feature_n = FeatureBuf_195;
         Mult_Buf[97].Weight_n = Wgt_1_195;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     end
    12:begin
     nxt_state = 13;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_196;
         Mult_Buf[0].Weight_n = Wgt_1_196;
         Mult_Buf[1].Feature_n = FeatureBuf_197;
         Mult_Buf[1].Weight_n = Wgt_1_197;
         Mult_Buf[2].Feature_n = FeatureBuf_198;
         Mult_Buf[2].Weight_n = Wgt_1_198;
         Mult_Buf[3].Feature_n = FeatureBuf_199;
         Mult_Buf[3].Weight_n = Wgt_1_199;
         Mult_Buf[4].Feature_n = FeatureBuf_200;
         Mult_Buf[4].Weight_n = Wgt_1_200;
         Mult_Buf[5].Feature_n = FeatureBuf_201;
         Mult_Buf[5].Weight_n = Wgt_1_201;
         Mult_Buf[6].Feature_n = FeatureBuf_202;
         Mult_Buf[6].Weight_n = Wgt_1_202;
         Mult_Buf[7].Feature_n = FeatureBuf_203;
         Mult_Buf[7].Weight_n = Wgt_1_203;
         Mult_Buf[8].Feature_n = FeatureBuf_204;
         Mult_Buf[8].Weight_n = Wgt_1_204;
         Mult_Buf[9].Feature_n = FeatureBuf_205;
         Mult_Buf[9].Weight_n = Wgt_1_205;
         Mult_Buf[10].Feature_n = FeatureBuf_206;
         Mult_Buf[10].Weight_n = Wgt_1_206;
         Mult_Buf[11].Feature_n = FeatureBuf_207;
         Mult_Buf[11].Weight_n = Wgt_1_207;
         Mult_Buf[12].Feature_n = FeatureBuf_208;
         Mult_Buf[12].Weight_n = Wgt_1_208;
         Mult_Buf[13].Feature_n = FeatureBuf_209;
         Mult_Buf[13].Weight_n = Wgt_1_209;
         Mult_Buf[14].Feature_n = FeatureBuf_210;
         Mult_Buf[14].Weight_n = Wgt_1_210;
         Mult_Buf[15].Feature_n = FeatureBuf_211;
         Mult_Buf[15].Weight_n = Wgt_1_211;
         Mult_Buf[16].Feature_n = FeatureBuf_212;
         Mult_Buf[16].Weight_n = Wgt_1_212;
         Mult_Buf[17].Feature_n = FeatureBuf_213;
         Mult_Buf[17].Weight_n = Wgt_1_213;
         Mult_Buf[18].Feature_n = FeatureBuf_214;
         Mult_Buf[18].Weight_n = Wgt_1_214;
         Mult_Buf[19].Feature_n = FeatureBuf_215;
         Mult_Buf[19].Weight_n = Wgt_1_215;
         Mult_Buf[20].Feature_n = FeatureBuf_216;
         Mult_Buf[20].Weight_n = Wgt_1_216;
         Mult_Buf[21].Feature_n = FeatureBuf_217;
         Mult_Buf[21].Weight_n = Wgt_1_217;
         Mult_Buf[22].Feature_n = FeatureBuf_218;
         Mult_Buf[22].Weight_n = Wgt_1_218;
         Mult_Buf[23].Feature_n = FeatureBuf_219;
         Mult_Buf[23].Weight_n = Wgt_1_219;
         Mult_Buf[24].Feature_n = FeatureBuf_220;
         Mult_Buf[24].Weight_n = Wgt_1_220;
         Mult_Buf[25].Feature_n = FeatureBuf_221;
         Mult_Buf[25].Weight_n = Wgt_1_221;
         Mult_Buf[26].Feature_n = FeatureBuf_222;
         Mult_Buf[26].Weight_n = Wgt_1_222;
         Mult_Buf[27].Feature_n = FeatureBuf_223;
         Mult_Buf[27].Weight_n = Wgt_1_223;
         Mult_Buf[28].Feature_n = FeatureBuf_224;
         Mult_Buf[28].Weight_n = Wgt_1_224;
         Mult_Buf[29].Feature_n = FeatureBuf_225;
         Mult_Buf[29].Weight_n = Wgt_1_225;
         Mult_Buf[30].Feature_n = FeatureBuf_226;
         Mult_Buf[30].Weight_n = Wgt_1_226;
         Mult_Buf[31].Feature_n = FeatureBuf_227;
         Mult_Buf[31].Weight_n = Wgt_1_227;
         Mult_Buf[32].Feature_n = FeatureBuf_228;
         Mult_Buf[32].Weight_n = Wgt_1_228;
         Mult_Buf[33].Feature_n = FeatureBuf_229;
         Mult_Buf[33].Weight_n = Wgt_1_229;
         Mult_Buf[34].Feature_n = FeatureBuf_230;
         Mult_Buf[34].Weight_n = Wgt_1_230;
         Mult_Buf[35].Feature_n = FeatureBuf_231;
         Mult_Buf[35].Weight_n = Wgt_1_231;
         Mult_Buf[36].Feature_n = FeatureBuf_232;
         Mult_Buf[36].Weight_n = Wgt_1_232;
         Mult_Buf[37].Feature_n = FeatureBuf_233;
         Mult_Buf[37].Weight_n = Wgt_1_233;
         Mult_Buf[38].Feature_n = FeatureBuf_234;
         Mult_Buf[38].Weight_n = Wgt_1_234;
         Mult_Buf[39].Feature_n = FeatureBuf_235;
         Mult_Buf[39].Weight_n = Wgt_1_235;
         Mult_Buf[40].Feature_n = FeatureBuf_236;
         Mult_Buf[40].Weight_n = Wgt_1_236;
         Mult_Buf[41].Feature_n = FeatureBuf_237;
         Mult_Buf[41].Weight_n = Wgt_1_237;
         Mult_Buf[42].Feature_n = FeatureBuf_238;
         Mult_Buf[42].Weight_n = Wgt_1_238;
         Mult_Buf[43].Feature_n = FeatureBuf_239;
         Mult_Buf[43].Weight_n = Wgt_1_239;
         Mult_Buf[44].Feature_n = FeatureBuf_240;
         Mult_Buf[44].Weight_n = Wgt_1_240;
         Mult_Buf[45].Feature_n = FeatureBuf_241;
         Mult_Buf[45].Weight_n = Wgt_1_241;
         Mult_Buf[46].Feature_n = FeatureBuf_242;
         Mult_Buf[46].Weight_n = Wgt_1_242;
         Mult_Buf[47].Feature_n = FeatureBuf_243;
         Mult_Buf[47].Weight_n = Wgt_1_243;
         Mult_Buf[48].Feature_n = FeatureBuf_244;
         Mult_Buf[48].Weight_n = Wgt_1_244;
         Mult_Buf[49].Feature_n = FeatureBuf_245;
         Mult_Buf[49].Weight_n = Wgt_1_245;
         Mult_Buf[50].Feature_n = FeatureBuf_246;
         Mult_Buf[50].Weight_n = Wgt_1_246;
         Mult_Buf[51].Feature_n = FeatureBuf_247;
         Mult_Buf[51].Weight_n = Wgt_1_247;
         Mult_Buf[52].Feature_n = FeatureBuf_248;
         Mult_Buf[52].Weight_n = Wgt_1_248;
         Mult_Buf[53].Feature_n = FeatureBuf_249;
         Mult_Buf[53].Weight_n = Wgt_1_249;
         Mult_Buf[54].Feature_n = FeatureBuf_250;
         Mult_Buf[54].Weight_n = Wgt_1_250;
         Mult_Buf[55].Feature_n = FeatureBuf_251;
         Mult_Buf[55].Weight_n = Wgt_1_251;
         Mult_Buf[56].Feature_n = FeatureBuf_252;
         Mult_Buf[56].Weight_n = Wgt_1_252;
         Mult_Buf[57].Feature_n = FeatureBuf_253;
         Mult_Buf[57].Weight_n = Wgt_1_253;
         Mult_Buf[58].Feature_n = FeatureBuf_254;
         Mult_Buf[58].Weight_n = Wgt_1_254;
         Mult_Buf[59].Feature_n = FeatureBuf_255;
         Mult_Buf[59].Weight_n = Wgt_1_255;
         Mult_Buf[60].Feature_n = FeatureBuf_256;
         Mult_Buf[60].Weight_n = Wgt_1_256;
         Mult_Buf[61].Feature_n = FeatureBuf_257;
         Mult_Buf[61].Weight_n = Wgt_1_257;
         Mult_Buf[62].Feature_n = FeatureBuf_258;
         Mult_Buf[62].Weight_n = Wgt_1_258;
         Mult_Buf[63].Feature_n = FeatureBuf_259;
         Mult_Buf[63].Weight_n = Wgt_1_259;
         Mult_Buf[64].Feature_n = FeatureBuf_260;
         Mult_Buf[64].Weight_n = Wgt_1_260;
         Mult_Buf[65].Feature_n = FeatureBuf_261;
         Mult_Buf[65].Weight_n = Wgt_1_261;
         Mult_Buf[66].Feature_n = FeatureBuf_262;
         Mult_Buf[66].Weight_n = Wgt_1_262;
         Mult_Buf[67].Feature_n = FeatureBuf_263;
         Mult_Buf[67].Weight_n = Wgt_1_263;
         Mult_Buf[68].Feature_n = FeatureBuf_264;
         Mult_Buf[68].Weight_n = Wgt_1_264;
         Mult_Buf[69].Feature_n = FeatureBuf_265;
         Mult_Buf[69].Weight_n = Wgt_1_265;
         Mult_Buf[70].Feature_n = FeatureBuf_266;
         Mult_Buf[70].Weight_n = Wgt_1_266;
         Mult_Buf[71].Feature_n = FeatureBuf_267;
         Mult_Buf[71].Weight_n = Wgt_1_267;
         Mult_Buf[72].Feature_n = FeatureBuf_268;
         Mult_Buf[72].Weight_n = Wgt_1_268;
         Mult_Buf[73].Feature_n = FeatureBuf_269;
         Mult_Buf[73].Weight_n = Wgt_1_269;
         Mult_Buf[74].Feature_n = FeatureBuf_270;
         Mult_Buf[74].Weight_n = Wgt_1_270;
         Mult_Buf[75].Feature_n = FeatureBuf_271;
         Mult_Buf[75].Weight_n = Wgt_1_271;
         Mult_Buf[76].Feature_n = FeatureBuf_272;
         Mult_Buf[76].Weight_n = Wgt_1_272;
         Mult_Buf[77].Feature_n = FeatureBuf_273;
         Mult_Buf[77].Weight_n = Wgt_1_273;
         Mult_Buf[78].Feature_n = FeatureBuf_274;
         Mult_Buf[78].Weight_n = Wgt_1_274;
         Mult_Buf[79].Feature_n = FeatureBuf_275;
         Mult_Buf[79].Weight_n = Wgt_1_275;
         Mult_Buf[80].Feature_n = FeatureBuf_276;
         Mult_Buf[80].Weight_n = Wgt_1_276;
         Mult_Buf[81].Feature_n = FeatureBuf_277;
         Mult_Buf[81].Weight_n = Wgt_1_277;
         Mult_Buf[82].Feature_n = FeatureBuf_278;
         Mult_Buf[82].Weight_n = Wgt_1_278;
         Mult_Buf[83].Feature_n = FeatureBuf_279;
         Mult_Buf[83].Weight_n = Wgt_1_279;
         Mult_Buf[84].Feature_n = FeatureBuf_280;
         Mult_Buf[84].Weight_n = Wgt_1_280;
         Mult_Buf[85].Feature_n = FeatureBuf_281;
         Mult_Buf[85].Weight_n = Wgt_1_281;
         Mult_Buf[86].Feature_n = FeatureBuf_282;
         Mult_Buf[86].Weight_n = Wgt_1_282;
         Mult_Buf[87].Feature_n = FeatureBuf_283;
         Mult_Buf[87].Weight_n = Wgt_1_283;
         Mult_Buf[88].Feature_n = FeatureBuf_284;
         Mult_Buf[88].Weight_n = Wgt_1_284;
         Mult_Buf[89].Feature_n = FeatureBuf_285;
         Mult_Buf[89].Weight_n = Wgt_1_285;
         Mult_Buf[90].Feature_n = FeatureBuf_286;
         Mult_Buf[90].Weight_n = Wgt_1_286;
         Mult_Buf[91].Feature_n = FeatureBuf_287;
         Mult_Buf[91].Weight_n = Wgt_1_287;
         Mult_Buf[92].Feature_n = FeatureBuf_288;
         Mult_Buf[92].Weight_n = Wgt_1_288;
         Mult_Buf[93].Feature_n = FeatureBuf_289;
         Mult_Buf[93].Weight_n = Wgt_1_289;
         Mult_Buf[94].Feature_n = FeatureBuf_290;
         Mult_Buf[94].Weight_n = Wgt_1_290;
         Mult_Buf[95].Feature_n = FeatureBuf_291;
         Mult_Buf[95].Weight_n = Wgt_1_291;
         Mult_Buf[96].Feature_n = FeatureBuf_292;
         Mult_Buf[96].Weight_n = Wgt_1_292;
         Mult_Buf[97].Feature_n = FeatureBuf_293;
         Mult_Buf[97].Weight_n = Wgt_1_293;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     end
    13:begin
     nxt_state = 14;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_294;
         Mult_Buf[0].Weight_n = Wgt_1_294;
         Mult_Buf[1].Feature_n = FeatureBuf_295;
         Mult_Buf[1].Weight_n = Wgt_1_295;
         Mult_Buf[2].Feature_n = FeatureBuf_296;
         Mult_Buf[2].Weight_n = Wgt_1_296;
         Mult_Buf[3].Feature_n = FeatureBuf_297;
         Mult_Buf[3].Weight_n = Wgt_1_297;
         Mult_Buf[4].Feature_n = FeatureBuf_298;
         Mult_Buf[4].Weight_n = Wgt_1_298;
         Mult_Buf[5].Feature_n = FeatureBuf_299;
         Mult_Buf[5].Weight_n = Wgt_1_299;
         Mult_Buf[6].Feature_n = FeatureBuf_300;
         Mult_Buf[6].Weight_n = Wgt_1_300;
         Mult_Buf[7].Feature_n = FeatureBuf_301;
         Mult_Buf[7].Weight_n = Wgt_1_301;
         Mult_Buf[8].Feature_n = FeatureBuf_302;
         Mult_Buf[8].Weight_n = Wgt_1_302;
         Mult_Buf[9].Feature_n = FeatureBuf_303;
         Mult_Buf[9].Weight_n = Wgt_1_303;
         Mult_Buf[10].Feature_n = FeatureBuf_304;
         Mult_Buf[10].Weight_n = Wgt_1_304;
         Mult_Buf[11].Feature_n = FeatureBuf_305;
         Mult_Buf[11].Weight_n = Wgt_1_305;
         Mult_Buf[12].Feature_n = FeatureBuf_306;
         Mult_Buf[12].Weight_n = Wgt_1_306;
         Mult_Buf[13].Feature_n = FeatureBuf_307;
         Mult_Buf[13].Weight_n = Wgt_1_307;
         Mult_Buf[14].Feature_n = FeatureBuf_308;
         Mult_Buf[14].Weight_n = Wgt_1_308;
         Mult_Buf[15].Feature_n = FeatureBuf_309;
         Mult_Buf[15].Weight_n = Wgt_1_309;
         Mult_Buf[16].Feature_n = FeatureBuf_310;
         Mult_Buf[16].Weight_n = Wgt_1_310;
         Mult_Buf[17].Feature_n = FeatureBuf_311;
         Mult_Buf[17].Weight_n = Wgt_1_311;
         Mult_Buf[18].Feature_n = FeatureBuf_312;
         Mult_Buf[18].Weight_n = Wgt_1_312;
         Mult_Buf[19].Feature_n = FeatureBuf_313;
         Mult_Buf[19].Weight_n = Wgt_1_313;
         Mult_Buf[20].Feature_n = FeatureBuf_314;
         Mult_Buf[20].Weight_n = Wgt_1_314;
         Mult_Buf[21].Feature_n = FeatureBuf_315;
         Mult_Buf[21].Weight_n = Wgt_1_315;
         Mult_Buf[22].Feature_n = FeatureBuf_316;
         Mult_Buf[22].Weight_n = Wgt_1_316;
         Mult_Buf[23].Feature_n = FeatureBuf_317;
         Mult_Buf[23].Weight_n = Wgt_1_317;
         Mult_Buf[24].Feature_n = FeatureBuf_318;
         Mult_Buf[24].Weight_n = Wgt_1_318;
         Mult_Buf[25].Feature_n = FeatureBuf_319;
         Mult_Buf[25].Weight_n = Wgt_1_319;
         Mult_Buf[26].Feature_n = FeatureBuf_320;
         Mult_Buf[26].Weight_n = Wgt_1_320;
         Mult_Buf[27].Feature_n = FeatureBuf_321;
         Mult_Buf[27].Weight_n = Wgt_1_321;
         Mult_Buf[28].Feature_n = FeatureBuf_322;
         Mult_Buf[28].Weight_n = Wgt_1_322;
         Mult_Buf[29].Feature_n = FeatureBuf_323;
         Mult_Buf[29].Weight_n = Wgt_1_323;
         Mult_Buf[30].Feature_n = FeatureBuf_324;
         Mult_Buf[30].Weight_n = Wgt_1_324;
         Mult_Buf[31].Feature_n = FeatureBuf_325;
         Mult_Buf[31].Weight_n = Wgt_1_325;
         Mult_Buf[32].Feature_n = FeatureBuf_326;
         Mult_Buf[32].Weight_n = Wgt_1_326;
         Mult_Buf[33].Feature_n = FeatureBuf_327;
         Mult_Buf[33].Weight_n = Wgt_1_327;
         Mult_Buf[34].Feature_n = FeatureBuf_328;
         Mult_Buf[34].Weight_n = Wgt_1_328;
         Mult_Buf[35].Feature_n = FeatureBuf_329;
         Mult_Buf[35].Weight_n = Wgt_1_329;
         Mult_Buf[36].Feature_n = FeatureBuf_330;
         Mult_Buf[36].Weight_n = Wgt_1_330;
         Mult_Buf[37].Feature_n = FeatureBuf_331;
         Mult_Buf[37].Weight_n = Wgt_1_331;
         Mult_Buf[38].Feature_n = FeatureBuf_332;
         Mult_Buf[38].Weight_n = Wgt_1_332;
         Mult_Buf[39].Feature_n = FeatureBuf_333;
         Mult_Buf[39].Weight_n = Wgt_1_333;
         Mult_Buf[40].Feature_n = FeatureBuf_334;
         Mult_Buf[40].Weight_n = Wgt_1_334;
         Mult_Buf[41].Feature_n = FeatureBuf_335;
         Mult_Buf[41].Weight_n = Wgt_1_335;
         Mult_Buf[42].Feature_n = FeatureBuf_336;
         Mult_Buf[42].Weight_n = Wgt_1_336;
         Mult_Buf[43].Feature_n = FeatureBuf_337;
         Mult_Buf[43].Weight_n = Wgt_1_337;
         Mult_Buf[44].Feature_n = FeatureBuf_338;
         Mult_Buf[44].Weight_n = Wgt_1_338;
         Mult_Buf[45].Feature_n = FeatureBuf_339;
         Mult_Buf[45].Weight_n = Wgt_1_339;
         Mult_Buf[46].Feature_n = FeatureBuf_340;
         Mult_Buf[46].Weight_n = Wgt_1_340;
         Mult_Buf[47].Feature_n = FeatureBuf_341;
         Mult_Buf[47].Weight_n = Wgt_1_341;
         Mult_Buf[48].Feature_n = FeatureBuf_342;
         Mult_Buf[48].Weight_n = Wgt_1_342;
         Mult_Buf[49].Feature_n = FeatureBuf_343;
         Mult_Buf[49].Weight_n = Wgt_1_343;
         Mult_Buf[50].Feature_n = FeatureBuf_344;
         Mult_Buf[50].Weight_n = Wgt_1_344;
         Mult_Buf[51].Feature_n = FeatureBuf_345;
         Mult_Buf[51].Weight_n = Wgt_1_345;
         Mult_Buf[52].Feature_n = FeatureBuf_346;
         Mult_Buf[52].Weight_n = Wgt_1_346;
         Mult_Buf[53].Feature_n = FeatureBuf_347;
         Mult_Buf[53].Weight_n = Wgt_1_347;
         Mult_Buf[54].Feature_n = FeatureBuf_348;
         Mult_Buf[54].Weight_n = Wgt_1_348;
         Mult_Buf[55].Feature_n = FeatureBuf_349;
         Mult_Buf[55].Weight_n = Wgt_1_349;
         Mult_Buf[56].Feature_n = FeatureBuf_350;
         Mult_Buf[56].Weight_n = Wgt_1_350;
         Mult_Buf[57].Feature_n = FeatureBuf_351;
         Mult_Buf[57].Weight_n = Wgt_1_351;
         Mult_Buf[58].Feature_n = FeatureBuf_352;
         Mult_Buf[58].Weight_n = Wgt_1_352;
         Mult_Buf[59].Feature_n = FeatureBuf_353;
         Mult_Buf[59].Weight_n = Wgt_1_353;
         Mult_Buf[60].Feature_n = FeatureBuf_354;
         Mult_Buf[60].Weight_n = Wgt_1_354;
         Mult_Buf[61].Feature_n = FeatureBuf_355;
         Mult_Buf[61].Weight_n = Wgt_1_355;
         Mult_Buf[62].Feature_n = FeatureBuf_356;
         Mult_Buf[62].Weight_n = Wgt_1_356;
         Mult_Buf[63].Feature_n = FeatureBuf_357;
         Mult_Buf[63].Weight_n = Wgt_1_357;
         Mult_Buf[64].Feature_n = FeatureBuf_358;
         Mult_Buf[64].Weight_n = Wgt_1_358;
         Mult_Buf[65].Feature_n = FeatureBuf_359;
         Mult_Buf[65].Weight_n = Wgt_1_359;
         Mult_Buf[66].Feature_n = FeatureBuf_360;
         Mult_Buf[66].Weight_n = Wgt_1_360;
         Mult_Buf[67].Feature_n = FeatureBuf_361;
         Mult_Buf[67].Weight_n = Wgt_1_361;
         Mult_Buf[68].Feature_n = FeatureBuf_362;
         Mult_Buf[68].Weight_n = Wgt_1_362;
         Mult_Buf[69].Feature_n = FeatureBuf_363;
         Mult_Buf[69].Weight_n = Wgt_1_363;
         Mult_Buf[70].Feature_n = FeatureBuf_364;
         Mult_Buf[70].Weight_n = Wgt_1_364;
         Mult_Buf[71].Feature_n = FeatureBuf_365;
         Mult_Buf[71].Weight_n = Wgt_1_365;
         Mult_Buf[72].Feature_n = FeatureBuf_366;
         Mult_Buf[72].Weight_n = Wgt_1_366;
         Mult_Buf[73].Feature_n = FeatureBuf_367;
         Mult_Buf[73].Weight_n = Wgt_1_367;
         Mult_Buf[74].Feature_n = FeatureBuf_368;
         Mult_Buf[74].Weight_n = Wgt_1_368;
         Mult_Buf[75].Feature_n = FeatureBuf_369;
         Mult_Buf[75].Weight_n = Wgt_1_369;
         Mult_Buf[76].Feature_n = FeatureBuf_370;
         Mult_Buf[76].Weight_n = Wgt_1_370;
         Mult_Buf[77].Feature_n = FeatureBuf_371;
         Mult_Buf[77].Weight_n = Wgt_1_371;
         Mult_Buf[78].Feature_n = FeatureBuf_372;
         Mult_Buf[78].Weight_n = Wgt_1_372;
         Mult_Buf[79].Feature_n = FeatureBuf_373;
         Mult_Buf[79].Weight_n = Wgt_1_373;
         Mult_Buf[80].Feature_n = FeatureBuf_374;
         Mult_Buf[80].Weight_n = Wgt_1_374;
         Mult_Buf[81].Feature_n = FeatureBuf_375;
         Mult_Buf[81].Weight_n = Wgt_1_375;
         Mult_Buf[82].Feature_n = FeatureBuf_376;
         Mult_Buf[82].Weight_n = Wgt_1_376;
         Mult_Buf[83].Feature_n = FeatureBuf_377;
         Mult_Buf[83].Weight_n = Wgt_1_377;
         Mult_Buf[84].Feature_n = FeatureBuf_378;
         Mult_Buf[84].Weight_n = Wgt_1_378;
         Mult_Buf[85].Feature_n = FeatureBuf_379;
         Mult_Buf[85].Weight_n = Wgt_1_379;
         Mult_Buf[86].Feature_n = FeatureBuf_380;
         Mult_Buf[86].Weight_n = Wgt_1_380;
         Mult_Buf[87].Feature_n = FeatureBuf_381;
         Mult_Buf[87].Weight_n = Wgt_1_381;
         Mult_Buf[88].Feature_n = FeatureBuf_382;
         Mult_Buf[88].Weight_n = Wgt_1_382;
         Mult_Buf[89].Feature_n = FeatureBuf_383;
         Mult_Buf[89].Weight_n = Wgt_1_383;
         Mult_Buf[90].Feature_n = FeatureBuf_384;
         Mult_Buf[90].Weight_n = Wgt_1_384;
         Mult_Buf[91].Feature_n = FeatureBuf_385;
         Mult_Buf[91].Weight_n = Wgt_1_385;
         Mult_Buf[92].Feature_n = FeatureBuf_386;
         Mult_Buf[92].Weight_n = Wgt_1_386;
         Mult_Buf[93].Feature_n = FeatureBuf_387;
         Mult_Buf[93].Weight_n = Wgt_1_387;
         Mult_Buf[94].Feature_n = FeatureBuf_388;
         Mult_Buf[94].Weight_n = Wgt_1_388;
         Mult_Buf[95].Feature_n = FeatureBuf_389;
         Mult_Buf[95].Weight_n = Wgt_1_389;
         Mult_Buf[96].Feature_n = FeatureBuf_390;
         Mult_Buf[96].Weight_n = Wgt_1_390;
         Mult_Buf[97].Feature_n = FeatureBuf_391;
         Mult_Buf[97].Weight_n = Wgt_1_391;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     end
    14:begin
     nxt_state = 15;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_392;
         Mult_Buf[0].Weight_n = Wgt_1_392;
         Mult_Buf[1].Feature_n = FeatureBuf_393;
         Mult_Buf[1].Weight_n = Wgt_1_393;
         Mult_Buf[2].Feature_n = FeatureBuf_394;
         Mult_Buf[2].Weight_n = Wgt_1_394;
         Mult_Buf[3].Feature_n = FeatureBuf_395;
         Mult_Buf[3].Weight_n = Wgt_1_395;
         Mult_Buf[4].Feature_n = FeatureBuf_396;
         Mult_Buf[4].Weight_n = Wgt_1_396;
         Mult_Buf[5].Feature_n = FeatureBuf_397;
         Mult_Buf[5].Weight_n = Wgt_1_397;
         Mult_Buf[6].Feature_n = FeatureBuf_398;
         Mult_Buf[6].Weight_n = Wgt_1_398;
         Mult_Buf[7].Feature_n = FeatureBuf_399;
         Mult_Buf[7].Weight_n = Wgt_1_399;
         Mult_Buf[8].Feature_n = FeatureBuf_400;
         Mult_Buf[8].Weight_n = Wgt_1_400;
         Mult_Buf[9].Feature_n = FeatureBuf_401;
         Mult_Buf[9].Weight_n = Wgt_1_401;
         Mult_Buf[10].Feature_n = FeatureBuf_402;
         Mult_Buf[10].Weight_n = Wgt_1_402;
         Mult_Buf[11].Feature_n = FeatureBuf_403;
         Mult_Buf[11].Weight_n = Wgt_1_403;
         Mult_Buf[12].Feature_n = FeatureBuf_404;
         Mult_Buf[12].Weight_n = Wgt_1_404;
         Mult_Buf[13].Feature_n = FeatureBuf_405;
         Mult_Buf[13].Weight_n = Wgt_1_405;
         Mult_Buf[14].Feature_n = FeatureBuf_406;
         Mult_Buf[14].Weight_n = Wgt_1_406;
         Mult_Buf[15].Feature_n = FeatureBuf_407;
         Mult_Buf[15].Weight_n = Wgt_1_407;
         Mult_Buf[16].Feature_n = FeatureBuf_408;
         Mult_Buf[16].Weight_n = Wgt_1_408;
         Mult_Buf[17].Feature_n = FeatureBuf_409;
         Mult_Buf[17].Weight_n = Wgt_1_409;
         Mult_Buf[18].Feature_n = FeatureBuf_410;
         Mult_Buf[18].Weight_n = Wgt_1_410;
         Mult_Buf[19].Feature_n = FeatureBuf_411;
         Mult_Buf[19].Weight_n = Wgt_1_411;
         Mult_Buf[20].Feature_n = FeatureBuf_412;
         Mult_Buf[20].Weight_n = Wgt_1_412;
         Mult_Buf[21].Feature_n = FeatureBuf_413;
         Mult_Buf[21].Weight_n = Wgt_1_413;
         Mult_Buf[22].Feature_n = FeatureBuf_414;
         Mult_Buf[22].Weight_n = Wgt_1_414;
         Mult_Buf[23].Feature_n = FeatureBuf_415;
         Mult_Buf[23].Weight_n = Wgt_1_415;
         Mult_Buf[24].Feature_n = FeatureBuf_416;
         Mult_Buf[24].Weight_n = Wgt_1_416;
         Mult_Buf[25].Feature_n = FeatureBuf_417;
         Mult_Buf[25].Weight_n = Wgt_1_417;
         Mult_Buf[26].Feature_n = FeatureBuf_418;
         Mult_Buf[26].Weight_n = Wgt_1_418;
         Mult_Buf[27].Feature_n = FeatureBuf_419;
         Mult_Buf[27].Weight_n = Wgt_1_419;
         Mult_Buf[28].Feature_n = FeatureBuf_420;
         Mult_Buf[28].Weight_n = Wgt_1_420;
         Mult_Buf[29].Feature_n = FeatureBuf_421;
         Mult_Buf[29].Weight_n = Wgt_1_421;
         Mult_Buf[30].Feature_n = FeatureBuf_422;
         Mult_Buf[30].Weight_n = Wgt_1_422;
         Mult_Buf[31].Feature_n = FeatureBuf_423;
         Mult_Buf[31].Weight_n = Wgt_1_423;
         Mult_Buf[32].Feature_n = FeatureBuf_424;
         Mult_Buf[32].Weight_n = Wgt_1_424;
         Mult_Buf[33].Feature_n = FeatureBuf_425;
         Mult_Buf[33].Weight_n = Wgt_1_425;
         Mult_Buf[34].Feature_n = FeatureBuf_426;
         Mult_Buf[34].Weight_n = Wgt_1_426;
         Mult_Buf[35].Feature_n = FeatureBuf_427;
         Mult_Buf[35].Weight_n = Wgt_1_427;
         Mult_Buf[36].Feature_n = FeatureBuf_428;
         Mult_Buf[36].Weight_n = Wgt_1_428;
         Mult_Buf[37].Feature_n = FeatureBuf_429;
         Mult_Buf[37].Weight_n = Wgt_1_429;
         Mult_Buf[38].Feature_n = FeatureBuf_430;
         Mult_Buf[38].Weight_n = Wgt_1_430;
         Mult_Buf[39].Feature_n = FeatureBuf_431;
         Mult_Buf[39].Weight_n = Wgt_1_431;
         Mult_Buf[40].Feature_n = FeatureBuf_432;
         Mult_Buf[40].Weight_n = Wgt_1_432;
         Mult_Buf[41].Feature_n = FeatureBuf_433;
         Mult_Buf[41].Weight_n = Wgt_1_433;
         Mult_Buf[42].Feature_n = FeatureBuf_434;
         Mult_Buf[42].Weight_n = Wgt_1_434;
         Mult_Buf[43].Feature_n = FeatureBuf_435;
         Mult_Buf[43].Weight_n = Wgt_1_435;
         Mult_Buf[44].Feature_n = FeatureBuf_436;
         Mult_Buf[44].Weight_n = Wgt_1_436;
         Mult_Buf[45].Feature_n = FeatureBuf_437;
         Mult_Buf[45].Weight_n = Wgt_1_437;
         Mult_Buf[46].Feature_n = FeatureBuf_438;
         Mult_Buf[46].Weight_n = Wgt_1_438;
         Mult_Buf[47].Feature_n = FeatureBuf_439;
         Mult_Buf[47].Weight_n = Wgt_1_439;
         Mult_Buf[48].Feature_n = FeatureBuf_440;
         Mult_Buf[48].Weight_n = Wgt_1_440;
         Mult_Buf[49].Feature_n = FeatureBuf_441;
         Mult_Buf[49].Weight_n = Wgt_1_441;
         Mult_Buf[50].Feature_n = FeatureBuf_442;
         Mult_Buf[50].Weight_n = Wgt_1_442;
         Mult_Buf[51].Feature_n = FeatureBuf_443;
         Mult_Buf[51].Weight_n = Wgt_1_443;
         Mult_Buf[52].Feature_n = FeatureBuf_444;
         Mult_Buf[52].Weight_n = Wgt_1_444;
         Mult_Buf[53].Feature_n = FeatureBuf_445;
         Mult_Buf[53].Weight_n = Wgt_1_445;
         Mult_Buf[54].Feature_n = FeatureBuf_446;
         Mult_Buf[54].Weight_n = Wgt_1_446;
         Mult_Buf[55].Feature_n = FeatureBuf_447;
         Mult_Buf[55].Weight_n = Wgt_1_447;
         Mult_Buf[56].Feature_n = FeatureBuf_448;
         Mult_Buf[56].Weight_n = Wgt_1_448;
         Mult_Buf[57].Feature_n = FeatureBuf_449;
         Mult_Buf[57].Weight_n = Wgt_1_449;
         Mult_Buf[58].Feature_n = FeatureBuf_450;
         Mult_Buf[58].Weight_n = Wgt_1_450;
         Mult_Buf[59].Feature_n = FeatureBuf_451;
         Mult_Buf[59].Weight_n = Wgt_1_451;
         Mult_Buf[60].Feature_n = FeatureBuf_452;
         Mult_Buf[60].Weight_n = Wgt_1_452;
         Mult_Buf[61].Feature_n = FeatureBuf_453;
         Mult_Buf[61].Weight_n = Wgt_1_453;
         Mult_Buf[62].Feature_n = FeatureBuf_454;
         Mult_Buf[62].Weight_n = Wgt_1_454;
         Mult_Buf[63].Feature_n = FeatureBuf_455;
         Mult_Buf[63].Weight_n = Wgt_1_455;
         Mult_Buf[64].Feature_n = FeatureBuf_456;
         Mult_Buf[64].Weight_n = Wgt_1_456;
         Mult_Buf[65].Feature_n = FeatureBuf_457;
         Mult_Buf[65].Weight_n = Wgt_1_457;
         Mult_Buf[66].Feature_n = FeatureBuf_458;
         Mult_Buf[66].Weight_n = Wgt_1_458;
         Mult_Buf[67].Feature_n = FeatureBuf_459;
         Mult_Buf[67].Weight_n = Wgt_1_459;
         Mult_Buf[68].Feature_n = FeatureBuf_460;
         Mult_Buf[68].Weight_n = Wgt_1_460;
         Mult_Buf[69].Feature_n = FeatureBuf_461;
         Mult_Buf[69].Weight_n = Wgt_1_461;
         Mult_Buf[70].Feature_n = FeatureBuf_462;
         Mult_Buf[70].Weight_n = Wgt_1_462;
         Mult_Buf[71].Feature_n = FeatureBuf_463;
         Mult_Buf[71].Weight_n = Wgt_1_463;
         Mult_Buf[72].Feature_n = FeatureBuf_464;
         Mult_Buf[72].Weight_n = Wgt_1_464;
         Mult_Buf[73].Feature_n = FeatureBuf_465;
         Mult_Buf[73].Weight_n = Wgt_1_465;
         Mult_Buf[74].Feature_n = FeatureBuf_466;
         Mult_Buf[74].Weight_n = Wgt_1_466;
         Mult_Buf[75].Feature_n = FeatureBuf_467;
         Mult_Buf[75].Weight_n = Wgt_1_467;
         Mult_Buf[76].Feature_n = FeatureBuf_468;
         Mult_Buf[76].Weight_n = Wgt_1_468;
         Mult_Buf[77].Feature_n = FeatureBuf_469;
         Mult_Buf[77].Weight_n = Wgt_1_469;
         Mult_Buf[78].Feature_n = FeatureBuf_470;
         Mult_Buf[78].Weight_n = Wgt_1_470;
         Mult_Buf[79].Feature_n = FeatureBuf_471;
         Mult_Buf[79].Weight_n = Wgt_1_471;
         Mult_Buf[80].Feature_n = FeatureBuf_472;
         Mult_Buf[80].Weight_n = Wgt_1_472;
         Mult_Buf[81].Feature_n = FeatureBuf_473;
         Mult_Buf[81].Weight_n = Wgt_1_473;
         Mult_Buf[82].Feature_n = FeatureBuf_474;
         Mult_Buf[82].Weight_n = Wgt_1_474;
         Mult_Buf[83].Feature_n = FeatureBuf_475;
         Mult_Buf[83].Weight_n = Wgt_1_475;
         Mult_Buf[84].Feature_n = FeatureBuf_476;
         Mult_Buf[84].Weight_n = Wgt_1_476;
         Mult_Buf[85].Feature_n = FeatureBuf_477;
         Mult_Buf[85].Weight_n = Wgt_1_477;
         Mult_Buf[86].Feature_n = FeatureBuf_478;
         Mult_Buf[86].Weight_n = Wgt_1_478;
         Mult_Buf[87].Feature_n = FeatureBuf_479;
         Mult_Buf[87].Weight_n = Wgt_1_479;
         Mult_Buf[88].Feature_n = FeatureBuf_480;
         Mult_Buf[88].Weight_n = Wgt_1_480;
         Mult_Buf[89].Feature_n = FeatureBuf_481;
         Mult_Buf[89].Weight_n = Wgt_1_481;
         Mult_Buf[90].Feature_n = FeatureBuf_482;
         Mult_Buf[90].Weight_n = Wgt_1_482;
         Mult_Buf[91].Feature_n = FeatureBuf_483;
         Mult_Buf[91].Weight_n = Wgt_1_483;
         Mult_Buf[92].Feature_n = FeatureBuf_484;
         Mult_Buf[92].Weight_n = Wgt_1_484;
         Mult_Buf[93].Feature_n = FeatureBuf_485;
         Mult_Buf[93].Weight_n = Wgt_1_485;
         Mult_Buf[94].Feature_n = FeatureBuf_486;
         Mult_Buf[94].Weight_n = Wgt_1_486;
         Mult_Buf[95].Feature_n = FeatureBuf_487;
         Mult_Buf[95].Weight_n = Wgt_1_487;
         Mult_Buf[96].Feature_n = FeatureBuf_488;
         Mult_Buf[96].Weight_n = Wgt_1_488;
         Mult_Buf[97].Feature_n = FeatureBuf_489;
         Mult_Buf[97].Weight_n = Wgt_1_489;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     end
    15:begin
     nxt_state = 16;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_490;
         Mult_Buf[0].Weight_n = Wgt_1_490;
         Mult_Buf[1].Feature_n = FeatureBuf_491;
         Mult_Buf[1].Weight_n = Wgt_1_491;
         Mult_Buf[2].Feature_n = FeatureBuf_492;
         Mult_Buf[2].Weight_n = Wgt_1_492;
         Mult_Buf[3].Feature_n = FeatureBuf_493;
         Mult_Buf[3].Weight_n = Wgt_1_493;
         Mult_Buf[4].Feature_n = FeatureBuf_494;
         Mult_Buf[4].Weight_n = Wgt_1_494;
         Mult_Buf[5].Feature_n = FeatureBuf_495;
         Mult_Buf[5].Weight_n = Wgt_1_495;
         Mult_Buf[6].Feature_n = FeatureBuf_496;
         Mult_Buf[6].Weight_n = Wgt_1_496;
         Mult_Buf[7].Feature_n = FeatureBuf_497;
         Mult_Buf[7].Weight_n = Wgt_1_497;
         Mult_Buf[8].Feature_n = FeatureBuf_498;
         Mult_Buf[8].Weight_n = Wgt_1_498;
         Mult_Buf[9].Feature_n = FeatureBuf_499;
         Mult_Buf[9].Weight_n = Wgt_1_499;
         Mult_Buf[10].Feature_n = FeatureBuf_500;
         Mult_Buf[10].Weight_n = Wgt_1_500;
         Mult_Buf[11].Feature_n = FeatureBuf_501;
         Mult_Buf[11].Weight_n = Wgt_1_501;
         Mult_Buf[12].Feature_n = FeatureBuf_502;
         Mult_Buf[12].Weight_n = Wgt_1_502;
         Mult_Buf[13].Feature_n = FeatureBuf_503;
         Mult_Buf[13].Weight_n = Wgt_1_503;
         Mult_Buf[14].Feature_n = FeatureBuf_504;
         Mult_Buf[14].Weight_n = Wgt_1_504;
         Mult_Buf[15].Feature_n = FeatureBuf_505;
         Mult_Buf[15].Weight_n = Wgt_1_505;
         Mult_Buf[16].Feature_n = FeatureBuf_506;
         Mult_Buf[16].Weight_n = Wgt_1_506;
         Mult_Buf[17].Feature_n = FeatureBuf_507;
         Mult_Buf[17].Weight_n = Wgt_1_507;
         Mult_Buf[18].Feature_n = FeatureBuf_508;
         Mult_Buf[18].Weight_n = Wgt_1_508;
         Mult_Buf[19].Feature_n = FeatureBuf_509;
         Mult_Buf[19].Weight_n = Wgt_1_509;
         Mult_Buf[20].Feature_n = FeatureBuf_510;
         Mult_Buf[20].Weight_n = Wgt_1_510;
         Mult_Buf[21].Feature_n = FeatureBuf_511;
         Mult_Buf[21].Weight_n = Wgt_1_511;
         Mult_Buf[22].Feature_n = FeatureBuf_512;
         Mult_Buf[22].Weight_n = Wgt_1_512;
         Mult_Buf[23].Feature_n = FeatureBuf_513;
         Mult_Buf[23].Weight_n = Wgt_1_513;
         Mult_Buf[24].Feature_n = FeatureBuf_514;
         Mult_Buf[24].Weight_n = Wgt_1_514;
         Mult_Buf[25].Feature_n = FeatureBuf_515;
         Mult_Buf[25].Weight_n = Wgt_1_515;
         Mult_Buf[26].Feature_n = FeatureBuf_516;
         Mult_Buf[26].Weight_n = Wgt_1_516;
         Mult_Buf[27].Feature_n = FeatureBuf_517;
         Mult_Buf[27].Weight_n = Wgt_1_517;
         Mult_Buf[28].Feature_n = FeatureBuf_518;
         Mult_Buf[28].Weight_n = Wgt_1_518;
         Mult_Buf[29].Feature_n = FeatureBuf_519;
         Mult_Buf[29].Weight_n = Wgt_1_519;
         Mult_Buf[30].Feature_n = FeatureBuf_520;
         Mult_Buf[30].Weight_n = Wgt_1_520;
         Mult_Buf[31].Feature_n = FeatureBuf_521;
         Mult_Buf[31].Weight_n = Wgt_1_521;
         Mult_Buf[32].Feature_n = FeatureBuf_522;
         Mult_Buf[32].Weight_n = Wgt_1_522;
         Mult_Buf[33].Feature_n = FeatureBuf_523;
         Mult_Buf[33].Weight_n = Wgt_1_523;
         Mult_Buf[34].Feature_n = FeatureBuf_524;
         Mult_Buf[34].Weight_n = Wgt_1_524;
         Mult_Buf[35].Feature_n = FeatureBuf_525;
         Mult_Buf[35].Weight_n = Wgt_1_525;
         Mult_Buf[36].Feature_n = FeatureBuf_526;
         Mult_Buf[36].Weight_n = Wgt_1_526;
         Mult_Buf[37].Feature_n = FeatureBuf_527;
         Mult_Buf[37].Weight_n = Wgt_1_527;
         Mult_Buf[38].Feature_n = FeatureBuf_528;
         Mult_Buf[38].Weight_n = Wgt_1_528;
         Mult_Buf[39].Feature_n = FeatureBuf_529;
         Mult_Buf[39].Weight_n = Wgt_1_529;
         Mult_Buf[40].Feature_n = FeatureBuf_530;
         Mult_Buf[40].Weight_n = Wgt_1_530;
         Mult_Buf[41].Feature_n = FeatureBuf_531;
         Mult_Buf[41].Weight_n = Wgt_1_531;
         Mult_Buf[42].Feature_n = FeatureBuf_532;
         Mult_Buf[42].Weight_n = Wgt_1_532;
         Mult_Buf[43].Feature_n = FeatureBuf_533;
         Mult_Buf[43].Weight_n = Wgt_1_533;
         Mult_Buf[44].Feature_n = FeatureBuf_534;
         Mult_Buf[44].Weight_n = Wgt_1_534;
         Mult_Buf[45].Feature_n = FeatureBuf_535;
         Mult_Buf[45].Weight_n = Wgt_1_535;
         Mult_Buf[46].Feature_n = FeatureBuf_536;
         Mult_Buf[46].Weight_n = Wgt_1_536;
         Mult_Buf[47].Feature_n = FeatureBuf_537;
         Mult_Buf[47].Weight_n = Wgt_1_537;
         Mult_Buf[48].Feature_n = FeatureBuf_538;
         Mult_Buf[48].Weight_n = Wgt_1_538;
         Mult_Buf[49].Feature_n = FeatureBuf_539;
         Mult_Buf[49].Weight_n = Wgt_1_539;
         Mult_Buf[50].Feature_n = FeatureBuf_540;
         Mult_Buf[50].Weight_n = Wgt_1_540;
         Mult_Buf[51].Feature_n = FeatureBuf_541;
         Mult_Buf[51].Weight_n = Wgt_1_541;
         Mult_Buf[52].Feature_n = FeatureBuf_542;
         Mult_Buf[52].Weight_n = Wgt_1_542;
         Mult_Buf[53].Feature_n = FeatureBuf_543;
         Mult_Buf[53].Weight_n = Wgt_1_543;
         Mult_Buf[54].Feature_n = FeatureBuf_544;
         Mult_Buf[54].Weight_n = Wgt_1_544;
         Mult_Buf[55].Feature_n = FeatureBuf_545;
         Mult_Buf[55].Weight_n = Wgt_1_545;
         Mult_Buf[56].Feature_n = FeatureBuf_546;
         Mult_Buf[56].Weight_n = Wgt_1_546;
         Mult_Buf[57].Feature_n = FeatureBuf_547;
         Mult_Buf[57].Weight_n = Wgt_1_547;
         Mult_Buf[58].Feature_n = FeatureBuf_548;
         Mult_Buf[58].Weight_n = Wgt_1_548;
         Mult_Buf[59].Feature_n = FeatureBuf_549;
         Mult_Buf[59].Weight_n = Wgt_1_549;
         Mult_Buf[60].Feature_n = FeatureBuf_550;
         Mult_Buf[60].Weight_n = Wgt_1_550;
         Mult_Buf[61].Feature_n = FeatureBuf_551;
         Mult_Buf[61].Weight_n = Wgt_1_551;
         Mult_Buf[62].Feature_n = FeatureBuf_552;
         Mult_Buf[62].Weight_n = Wgt_1_552;
         Mult_Buf[63].Feature_n = FeatureBuf_553;
         Mult_Buf[63].Weight_n = Wgt_1_553;
         Mult_Buf[64].Feature_n = FeatureBuf_554;
         Mult_Buf[64].Weight_n = Wgt_1_554;
         Mult_Buf[65].Feature_n = FeatureBuf_555;
         Mult_Buf[65].Weight_n = Wgt_1_555;
         Mult_Buf[66].Feature_n = FeatureBuf_556;
         Mult_Buf[66].Weight_n = Wgt_1_556;
         Mult_Buf[67].Feature_n = FeatureBuf_557;
         Mult_Buf[67].Weight_n = Wgt_1_557;
         Mult_Buf[68].Feature_n = FeatureBuf_558;
         Mult_Buf[68].Weight_n = Wgt_1_558;
         Mult_Buf[69].Feature_n = FeatureBuf_559;
         Mult_Buf[69].Weight_n = Wgt_1_559;
         Mult_Buf[70].Feature_n = FeatureBuf_560;
         Mult_Buf[70].Weight_n = Wgt_1_560;
         Mult_Buf[71].Feature_n = FeatureBuf_561;
         Mult_Buf[71].Weight_n = Wgt_1_561;
         Mult_Buf[72].Feature_n = FeatureBuf_562;
         Mult_Buf[72].Weight_n = Wgt_1_562;
         Mult_Buf[73].Feature_n = FeatureBuf_563;
         Mult_Buf[73].Weight_n = Wgt_1_563;
         Mult_Buf[74].Feature_n = FeatureBuf_564;
         Mult_Buf[74].Weight_n = Wgt_1_564;
         Mult_Buf[75].Feature_n = FeatureBuf_565;
         Mult_Buf[75].Weight_n = Wgt_1_565;
         Mult_Buf[76].Feature_n = FeatureBuf_566;
         Mult_Buf[76].Weight_n = Wgt_1_566;
         Mult_Buf[77].Feature_n = FeatureBuf_567;
         Mult_Buf[77].Weight_n = Wgt_1_567;
         Mult_Buf[78].Feature_n = FeatureBuf_568;
         Mult_Buf[78].Weight_n = Wgt_1_568;
         Mult_Buf[79].Feature_n = FeatureBuf_569;
         Mult_Buf[79].Weight_n = Wgt_1_569;
         Mult_Buf[80].Feature_n = FeatureBuf_570;
         Mult_Buf[80].Weight_n = Wgt_1_570;
         Mult_Buf[81].Feature_n = FeatureBuf_571;
         Mult_Buf[81].Weight_n = Wgt_1_571;
         Mult_Buf[82].Feature_n = FeatureBuf_572;
         Mult_Buf[82].Weight_n = Wgt_1_572;
         Mult_Buf[83].Feature_n = FeatureBuf_573;
         Mult_Buf[83].Weight_n = Wgt_1_573;
         Mult_Buf[84].Feature_n = FeatureBuf_574;
         Mult_Buf[84].Weight_n = Wgt_1_574;
         Mult_Buf[85].Feature_n = FeatureBuf_575;
         Mult_Buf[85].Weight_n = Wgt_1_575;
         Mult_Buf[86].Feature_n = FeatureBuf_576;
         Mult_Buf[86].Weight_n = Wgt_1_576;
         Mult_Buf[87].Feature_n = FeatureBuf_577;
         Mult_Buf[87].Weight_n = Wgt_1_577;
         Mult_Buf[88].Feature_n = FeatureBuf_578;
         Mult_Buf[88].Weight_n = Wgt_1_578;
         Mult_Buf[89].Feature_n = FeatureBuf_579;
         Mult_Buf[89].Weight_n = Wgt_1_579;
         Mult_Buf[90].Feature_n = FeatureBuf_580;
         Mult_Buf[90].Weight_n = Wgt_1_580;
         Mult_Buf[91].Feature_n = FeatureBuf_581;
         Mult_Buf[91].Weight_n = Wgt_1_581;
         Mult_Buf[92].Feature_n = FeatureBuf_582;
         Mult_Buf[92].Weight_n = Wgt_1_582;
         Mult_Buf[93].Feature_n = FeatureBuf_583;
         Mult_Buf[93].Weight_n = Wgt_1_583;
         Mult_Buf[94].Feature_n = FeatureBuf_584;
         Mult_Buf[94].Weight_n = Wgt_1_584;
         Mult_Buf[95].Feature_n = FeatureBuf_585;
         Mult_Buf[95].Weight_n = Wgt_1_585;
         Mult_Buf[96].Feature_n = FeatureBuf_586;
         Mult_Buf[96].Weight_n = Wgt_1_586;
         Mult_Buf[97].Feature_n = FeatureBuf_587;
         Mult_Buf[97].Weight_n = Wgt_1_587;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     end
    16:begin
     nxt_state = 17;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_588;
         Mult_Buf[0].Weight_n = Wgt_1_588;
         Mult_Buf[1].Feature_n = FeatureBuf_589;
         Mult_Buf[1].Weight_n = Wgt_1_589;
         Mult_Buf[2].Feature_n = FeatureBuf_590;
         Mult_Buf[2].Weight_n = Wgt_1_590;
         Mult_Buf[3].Feature_n = FeatureBuf_591;
         Mult_Buf[3].Weight_n = Wgt_1_591;
         Mult_Buf[4].Feature_n = FeatureBuf_592;
         Mult_Buf[4].Weight_n = Wgt_1_592;
         Mult_Buf[5].Feature_n = FeatureBuf_593;
         Mult_Buf[5].Weight_n = Wgt_1_593;
         Mult_Buf[6].Feature_n = FeatureBuf_594;
         Mult_Buf[6].Weight_n = Wgt_1_594;
         Mult_Buf[7].Feature_n = FeatureBuf_595;
         Mult_Buf[7].Weight_n = Wgt_1_595;
         Mult_Buf[8].Feature_n = FeatureBuf_596;
         Mult_Buf[8].Weight_n = Wgt_1_596;
         Mult_Buf[9].Feature_n = FeatureBuf_597;
         Mult_Buf[9].Weight_n = Wgt_1_597;
         Mult_Buf[10].Feature_n = FeatureBuf_598;
         Mult_Buf[10].Weight_n = Wgt_1_598;
         Mult_Buf[11].Feature_n = FeatureBuf_599;
         Mult_Buf[11].Weight_n = Wgt_1_599;
         Mult_Buf[12].Feature_n = FeatureBuf_600;
         Mult_Buf[12].Weight_n = Wgt_1_600;
         Mult_Buf[13].Feature_n = FeatureBuf_601;
         Mult_Buf[13].Weight_n = Wgt_1_601;
         Mult_Buf[14].Feature_n = FeatureBuf_602;
         Mult_Buf[14].Weight_n = Wgt_1_602;
         Mult_Buf[15].Feature_n = FeatureBuf_603;
         Mult_Buf[15].Weight_n = Wgt_1_603;
         Mult_Buf[16].Feature_n = FeatureBuf_604;
         Mult_Buf[16].Weight_n = Wgt_1_604;
         Mult_Buf[17].Feature_n = FeatureBuf_605;
         Mult_Buf[17].Weight_n = Wgt_1_605;
         Mult_Buf[18].Feature_n = FeatureBuf_606;
         Mult_Buf[18].Weight_n = Wgt_1_606;
         Mult_Buf[19].Feature_n = FeatureBuf_607;
         Mult_Buf[19].Weight_n = Wgt_1_607;
         Mult_Buf[20].Feature_n = FeatureBuf_608;
         Mult_Buf[20].Weight_n = Wgt_1_608;
         Mult_Buf[21].Feature_n = FeatureBuf_609;
         Mult_Buf[21].Weight_n = Wgt_1_609;
         Mult_Buf[22].Feature_n = FeatureBuf_610;
         Mult_Buf[22].Weight_n = Wgt_1_610;
         Mult_Buf[23].Feature_n = FeatureBuf_611;
         Mult_Buf[23].Weight_n = Wgt_1_611;
         Mult_Buf[24].Feature_n = FeatureBuf_612;
         Mult_Buf[24].Weight_n = Wgt_1_612;
         Mult_Buf[25].Feature_n = FeatureBuf_613;
         Mult_Buf[25].Weight_n = Wgt_1_613;
         Mult_Buf[26].Feature_n = FeatureBuf_614;
         Mult_Buf[26].Weight_n = Wgt_1_614;
         Mult_Buf[27].Feature_n = FeatureBuf_615;
         Mult_Buf[27].Weight_n = Wgt_1_615;
         Mult_Buf[28].Feature_n = FeatureBuf_616;
         Mult_Buf[28].Weight_n = Wgt_1_616;
         Mult_Buf[29].Feature_n = FeatureBuf_617;
         Mult_Buf[29].Weight_n = Wgt_1_617;
         Mult_Buf[30].Feature_n = FeatureBuf_618;
         Mult_Buf[30].Weight_n = Wgt_1_618;
         Mult_Buf[31].Feature_n = FeatureBuf_619;
         Mult_Buf[31].Weight_n = Wgt_1_619;
         Mult_Buf[32].Feature_n = FeatureBuf_620;
         Mult_Buf[32].Weight_n = Wgt_1_620;
         Mult_Buf[33].Feature_n = FeatureBuf_621;
         Mult_Buf[33].Weight_n = Wgt_1_621;
         Mult_Buf[34].Feature_n = FeatureBuf_622;
         Mult_Buf[34].Weight_n = Wgt_1_622;
         Mult_Buf[35].Feature_n = FeatureBuf_623;
         Mult_Buf[35].Weight_n = Wgt_1_623;
         Mult_Buf[36].Feature_n = FeatureBuf_624;
         Mult_Buf[36].Weight_n = Wgt_1_624;
         Mult_Buf[37].Feature_n = FeatureBuf_625;
         Mult_Buf[37].Weight_n = Wgt_1_625;
         Mult_Buf[38].Feature_n = FeatureBuf_626;
         Mult_Buf[38].Weight_n = Wgt_1_626;
         Mult_Buf[39].Feature_n = FeatureBuf_627;
         Mult_Buf[39].Weight_n = Wgt_1_627;
         Mult_Buf[40].Feature_n = FeatureBuf_628;
         Mult_Buf[40].Weight_n = Wgt_1_628;
         Mult_Buf[41].Feature_n = FeatureBuf_629;
         Mult_Buf[41].Weight_n = Wgt_1_629;
         Mult_Buf[42].Feature_n = FeatureBuf_630;
         Mult_Buf[42].Weight_n = Wgt_1_630;
         Mult_Buf[43].Feature_n = FeatureBuf_631;
         Mult_Buf[43].Weight_n = Wgt_1_631;
         Mult_Buf[44].Feature_n = FeatureBuf_632;
         Mult_Buf[44].Weight_n = Wgt_1_632;
         Mult_Buf[45].Feature_n = FeatureBuf_633;
         Mult_Buf[45].Weight_n = Wgt_1_633;
         Mult_Buf[46].Feature_n = FeatureBuf_634;
         Mult_Buf[46].Weight_n = Wgt_1_634;
         Mult_Buf[47].Feature_n = FeatureBuf_635;
         Mult_Buf[47].Weight_n = Wgt_1_635;
         Mult_Buf[48].Feature_n = FeatureBuf_636;
         Mult_Buf[48].Weight_n = Wgt_1_636;
         Mult_Buf[49].Feature_n = FeatureBuf_637;
         Mult_Buf[49].Weight_n = Wgt_1_637;
         Mult_Buf[50].Feature_n = FeatureBuf_638;
         Mult_Buf[50].Weight_n = Wgt_1_638;
         Mult_Buf[51].Feature_n = FeatureBuf_639;
         Mult_Buf[51].Weight_n = Wgt_1_639;
         Mult_Buf[52].Feature_n = FeatureBuf_640;
         Mult_Buf[52].Weight_n = Wgt_1_640;
         Mult_Buf[53].Feature_n = FeatureBuf_641;
         Mult_Buf[53].Weight_n = Wgt_1_641;
         Mult_Buf[54].Feature_n = FeatureBuf_642;
         Mult_Buf[54].Weight_n = Wgt_1_642;
         Mult_Buf[55].Feature_n = FeatureBuf_643;
         Mult_Buf[55].Weight_n = Wgt_1_643;
         Mult_Buf[56].Feature_n = FeatureBuf_644;
         Mult_Buf[56].Weight_n = Wgt_1_644;
         Mult_Buf[57].Feature_n = FeatureBuf_645;
         Mult_Buf[57].Weight_n = Wgt_1_645;
         Mult_Buf[58].Feature_n = FeatureBuf_646;
         Mult_Buf[58].Weight_n = Wgt_1_646;
         Mult_Buf[59].Feature_n = FeatureBuf_647;
         Mult_Buf[59].Weight_n = Wgt_1_647;
         Mult_Buf[60].Feature_n = FeatureBuf_648;
         Mult_Buf[60].Weight_n = Wgt_1_648;
         Mult_Buf[61].Feature_n = FeatureBuf_649;
         Mult_Buf[61].Weight_n = Wgt_1_649;
         Mult_Buf[62].Feature_n = FeatureBuf_650;
         Mult_Buf[62].Weight_n = Wgt_1_650;
         Mult_Buf[63].Feature_n = FeatureBuf_651;
         Mult_Buf[63].Weight_n = Wgt_1_651;
         Mult_Buf[64].Feature_n = FeatureBuf_652;
         Mult_Buf[64].Weight_n = Wgt_1_652;
         Mult_Buf[65].Feature_n = FeatureBuf_653;
         Mult_Buf[65].Weight_n = Wgt_1_653;
         Mult_Buf[66].Feature_n = FeatureBuf_654;
         Mult_Buf[66].Weight_n = Wgt_1_654;
         Mult_Buf[67].Feature_n = FeatureBuf_655;
         Mult_Buf[67].Weight_n = Wgt_1_655;
         Mult_Buf[68].Feature_n = FeatureBuf_656;
         Mult_Buf[68].Weight_n = Wgt_1_656;
         Mult_Buf[69].Feature_n = FeatureBuf_657;
         Mult_Buf[69].Weight_n = Wgt_1_657;
         Mult_Buf[70].Feature_n = FeatureBuf_658;
         Mult_Buf[70].Weight_n = Wgt_1_658;
         Mult_Buf[71].Feature_n = FeatureBuf_659;
         Mult_Buf[71].Weight_n = Wgt_1_659;
         Mult_Buf[72].Feature_n = FeatureBuf_660;
         Mult_Buf[72].Weight_n = Wgt_1_660;
         Mult_Buf[73].Feature_n = FeatureBuf_661;
         Mult_Buf[73].Weight_n = Wgt_1_661;
         Mult_Buf[74].Feature_n = FeatureBuf_662;
         Mult_Buf[74].Weight_n = Wgt_1_662;
         Mult_Buf[75].Feature_n = FeatureBuf_663;
         Mult_Buf[75].Weight_n = Wgt_1_663;
         Mult_Buf[76].Feature_n = FeatureBuf_664;
         Mult_Buf[76].Weight_n = Wgt_1_664;
         Mult_Buf[77].Feature_n = FeatureBuf_665;
         Mult_Buf[77].Weight_n = Wgt_1_665;
         Mult_Buf[78].Feature_n = FeatureBuf_666;
         Mult_Buf[78].Weight_n = Wgt_1_666;
         Mult_Buf[79].Feature_n = FeatureBuf_667;
         Mult_Buf[79].Weight_n = Wgt_1_667;
         Mult_Buf[80].Feature_n = FeatureBuf_668;
         Mult_Buf[80].Weight_n = Wgt_1_668;
         Mult_Buf[81].Feature_n = FeatureBuf_669;
         Mult_Buf[81].Weight_n = Wgt_1_669;
         Mult_Buf[82].Feature_n = FeatureBuf_670;
         Mult_Buf[82].Weight_n = Wgt_1_670;
         Mult_Buf[83].Feature_n = FeatureBuf_671;
         Mult_Buf[83].Weight_n = Wgt_1_671;
         Mult_Buf[84].Feature_n = FeatureBuf_672;
         Mult_Buf[84].Weight_n = Wgt_1_672;
         Mult_Buf[85].Feature_n = FeatureBuf_673;
         Mult_Buf[85].Weight_n = Wgt_1_673;
         Mult_Buf[86].Feature_n = FeatureBuf_674;
         Mult_Buf[86].Weight_n = Wgt_1_674;
         Mult_Buf[87].Feature_n = FeatureBuf_675;
         Mult_Buf[87].Weight_n = Wgt_1_675;
         Mult_Buf[88].Feature_n = FeatureBuf_676;
         Mult_Buf[88].Weight_n = Wgt_1_676;
         Mult_Buf[89].Feature_n = FeatureBuf_677;
         Mult_Buf[89].Weight_n = Wgt_1_677;
         Mult_Buf[90].Feature_n = FeatureBuf_678;
         Mult_Buf[90].Weight_n = Wgt_1_678;
         Mult_Buf[91].Feature_n = FeatureBuf_679;
         Mult_Buf[91].Weight_n = Wgt_1_679;
         Mult_Buf[92].Feature_n = FeatureBuf_680;
         Mult_Buf[92].Weight_n = Wgt_1_680;
         Mult_Buf[93].Feature_n = FeatureBuf_681;
         Mult_Buf[93].Weight_n = Wgt_1_681;
         Mult_Buf[94].Feature_n = FeatureBuf_682;
         Mult_Buf[94].Weight_n = Wgt_1_682;
         Mult_Buf[95].Feature_n = FeatureBuf_683;
         Mult_Buf[95].Weight_n = Wgt_1_683;
         Mult_Buf[96].Feature_n = FeatureBuf_684;
         Mult_Buf[96].Weight_n = Wgt_1_684;
         Mult_Buf[97].Feature_n = FeatureBuf_685;
         Mult_Buf[97].Weight_n = Wgt_1_685;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     end
    17:begin
     nxt_state = 18;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_686;
         Mult_Buf[0].Weight_n = Wgt_1_686;
         Mult_Buf[1].Feature_n = FeatureBuf_687;
         Mult_Buf[1].Weight_n = Wgt_1_687;
         Mult_Buf[2].Feature_n = FeatureBuf_688;
         Mult_Buf[2].Weight_n = Wgt_1_688;
         Mult_Buf[3].Feature_n = FeatureBuf_689;
         Mult_Buf[3].Weight_n = Wgt_1_689;
         Mult_Buf[4].Feature_n = FeatureBuf_690;
         Mult_Buf[4].Weight_n = Wgt_1_690;
         Mult_Buf[5].Feature_n = FeatureBuf_691;
         Mult_Buf[5].Weight_n = Wgt_1_691;
         Mult_Buf[6].Feature_n = FeatureBuf_692;
         Mult_Buf[6].Weight_n = Wgt_1_692;
         Mult_Buf[7].Feature_n = FeatureBuf_693;
         Mult_Buf[7].Weight_n = Wgt_1_693;
         Mult_Buf[8].Feature_n = FeatureBuf_694;
         Mult_Buf[8].Weight_n = Wgt_1_694;
         Mult_Buf[9].Feature_n = FeatureBuf_695;
         Mult_Buf[9].Weight_n = Wgt_1_695;
         Mult_Buf[10].Feature_n = FeatureBuf_696;
         Mult_Buf[10].Weight_n = Wgt_1_696;
         Mult_Buf[11].Feature_n = FeatureBuf_697;
         Mult_Buf[11].Weight_n = Wgt_1_697;
         Mult_Buf[12].Feature_n = FeatureBuf_698;
         Mult_Buf[12].Weight_n = Wgt_1_698;
         Mult_Buf[13].Feature_n = FeatureBuf_699;
         Mult_Buf[13].Weight_n = Wgt_1_699;
         Mult_Buf[14].Feature_n = FeatureBuf_700;
         Mult_Buf[14].Weight_n = Wgt_1_700;
         Mult_Buf[15].Feature_n = FeatureBuf_701;
         Mult_Buf[15].Weight_n = Wgt_1_701;
         Mult_Buf[16].Feature_n = FeatureBuf_702;
         Mult_Buf[16].Weight_n = Wgt_1_702;
         Mult_Buf[17].Feature_n = FeatureBuf_703;
         Mult_Buf[17].Weight_n = Wgt_1_703;
         Mult_Buf[18].Feature_n = FeatureBuf_704;
         Mult_Buf[18].Weight_n = Wgt_1_704;
         Mult_Buf[19].Feature_n = FeatureBuf_705;
         Mult_Buf[19].Weight_n = Wgt_1_705;
         Mult_Buf[20].Feature_n = FeatureBuf_706;
         Mult_Buf[20].Weight_n = Wgt_1_706;
         Mult_Buf[21].Feature_n = FeatureBuf_707;
         Mult_Buf[21].Weight_n = Wgt_1_707;
         Mult_Buf[22].Feature_n = FeatureBuf_708;
         Mult_Buf[22].Weight_n = Wgt_1_708;
         Mult_Buf[23].Feature_n = FeatureBuf_709;
         Mult_Buf[23].Weight_n = Wgt_1_709;
         Mult_Buf[24].Feature_n = FeatureBuf_710;
         Mult_Buf[24].Weight_n = Wgt_1_710;
         Mult_Buf[25].Feature_n = FeatureBuf_711;
         Mult_Buf[25].Weight_n = Wgt_1_711;
         Mult_Buf[26].Feature_n = FeatureBuf_712;
         Mult_Buf[26].Weight_n = Wgt_1_712;
         Mult_Buf[27].Feature_n = FeatureBuf_713;
         Mult_Buf[27].Weight_n = Wgt_1_713;
         Mult_Buf[28].Feature_n = FeatureBuf_714;
         Mult_Buf[28].Weight_n = Wgt_1_714;
         Mult_Buf[29].Feature_n = FeatureBuf_715;
         Mult_Buf[29].Weight_n = Wgt_1_715;
         Mult_Buf[30].Feature_n = FeatureBuf_716;
         Mult_Buf[30].Weight_n = Wgt_1_716;
         Mult_Buf[31].Feature_n = FeatureBuf_717;
         Mult_Buf[31].Weight_n = Wgt_1_717;
         Mult_Buf[32].Feature_n = FeatureBuf_718;
         Mult_Buf[32].Weight_n = Wgt_1_718;
         Mult_Buf[33].Feature_n = FeatureBuf_719;
         Mult_Buf[33].Weight_n = Wgt_1_719;
         Mult_Buf[34].Feature_n = FeatureBuf_720;
         Mult_Buf[34].Weight_n = Wgt_1_720;
         Mult_Buf[35].Feature_n = FeatureBuf_721;
         Mult_Buf[35].Weight_n = Wgt_1_721;
         Mult_Buf[36].Feature_n = FeatureBuf_722;
         Mult_Buf[36].Weight_n = Wgt_1_722;
         Mult_Buf[37].Feature_n = FeatureBuf_723;
         Mult_Buf[37].Weight_n = Wgt_1_723;
         Mult_Buf[38].Feature_n = FeatureBuf_724;
         Mult_Buf[38].Weight_n = Wgt_1_724;
         Mult_Buf[39].Feature_n = FeatureBuf_725;
         Mult_Buf[39].Weight_n = Wgt_1_725;
         Mult_Buf[40].Feature_n = FeatureBuf_726;
         Mult_Buf[40].Weight_n = Wgt_1_726;
         Mult_Buf[41].Feature_n = FeatureBuf_727;
         Mult_Buf[41].Weight_n = Wgt_1_727;
         Mult_Buf[42].Feature_n = FeatureBuf_728;
         Mult_Buf[42].Weight_n = Wgt_1_728;
         Mult_Buf[43].Feature_n = FeatureBuf_729;
         Mult_Buf[43].Weight_n = Wgt_1_729;
         Mult_Buf[44].Feature_n = FeatureBuf_730;
         Mult_Buf[44].Weight_n = Wgt_1_730;
         Mult_Buf[45].Feature_n = FeatureBuf_731;
         Mult_Buf[45].Weight_n = Wgt_1_731;
         Mult_Buf[46].Feature_n = FeatureBuf_732;
         Mult_Buf[46].Weight_n = Wgt_1_732;
         Mult_Buf[47].Feature_n = FeatureBuf_733;
         Mult_Buf[47].Weight_n = Wgt_1_733;
         Mult_Buf[48].Feature_n = FeatureBuf_734;
         Mult_Buf[48].Weight_n = Wgt_1_734;
         Mult_Buf[49].Feature_n = FeatureBuf_735;
         Mult_Buf[49].Weight_n = Wgt_1_735;
         Mult_Buf[50].Feature_n = FeatureBuf_736;
         Mult_Buf[50].Weight_n = Wgt_1_736;
         Mult_Buf[51].Feature_n = FeatureBuf_737;
         Mult_Buf[51].Weight_n = Wgt_1_737;
         Mult_Buf[52].Feature_n = FeatureBuf_738;
         Mult_Buf[52].Weight_n = Wgt_1_738;
         Mult_Buf[53].Feature_n = FeatureBuf_739;
         Mult_Buf[53].Weight_n = Wgt_1_739;
         Mult_Buf[54].Feature_n = FeatureBuf_740;
         Mult_Buf[54].Weight_n = Wgt_1_740;
         Mult_Buf[55].Feature_n = FeatureBuf_741;
         Mult_Buf[55].Weight_n = Wgt_1_741;
         Mult_Buf[56].Feature_n = FeatureBuf_742;
         Mult_Buf[56].Weight_n = Wgt_1_742;
         Mult_Buf[57].Feature_n = FeatureBuf_743;
         Mult_Buf[57].Weight_n = Wgt_1_743;
         Mult_Buf[58].Feature_n = FeatureBuf_744;
         Mult_Buf[58].Weight_n = Wgt_1_744;
         Mult_Buf[59].Feature_n = FeatureBuf_745;
         Mult_Buf[59].Weight_n = Wgt_1_745;
         Mult_Buf[60].Feature_n = FeatureBuf_746;
         Mult_Buf[60].Weight_n = Wgt_1_746;
         Mult_Buf[61].Feature_n = FeatureBuf_747;
         Mult_Buf[61].Weight_n = Wgt_1_747;
         Mult_Buf[62].Feature_n = FeatureBuf_748;
         Mult_Buf[62].Weight_n = Wgt_1_748;
         Mult_Buf[63].Feature_n = FeatureBuf_749;
         Mult_Buf[63].Weight_n = Wgt_1_749;
         Mult_Buf[64].Feature_n = FeatureBuf_750;
         Mult_Buf[64].Weight_n = Wgt_1_750;
         Mult_Buf[65].Feature_n = FeatureBuf_751;
         Mult_Buf[65].Weight_n = Wgt_1_751;
         Mult_Buf[66].Feature_n = FeatureBuf_752;
         Mult_Buf[66].Weight_n = Wgt_1_752;
         Mult_Buf[67].Feature_n = FeatureBuf_753;
         Mult_Buf[67].Weight_n = Wgt_1_753;
         Mult_Buf[68].Feature_n = FeatureBuf_754;
         Mult_Buf[68].Weight_n = Wgt_1_754;
         Mult_Buf[69].Feature_n = FeatureBuf_755;
         Mult_Buf[69].Weight_n = Wgt_1_755;
         Mult_Buf[70].Feature_n = FeatureBuf_756;
         Mult_Buf[70].Weight_n = Wgt_1_756;
         Mult_Buf[71].Feature_n = FeatureBuf_757;
         Mult_Buf[71].Weight_n = Wgt_1_757;
         Mult_Buf[72].Feature_n = FeatureBuf_758;
         Mult_Buf[72].Weight_n = Wgt_1_758;
         Mult_Buf[73].Feature_n = FeatureBuf_759;
         Mult_Buf[73].Weight_n = Wgt_1_759;
         Mult_Buf[74].Feature_n = FeatureBuf_760;
         Mult_Buf[74].Weight_n = Wgt_1_760;
         Mult_Buf[75].Feature_n = FeatureBuf_761;
         Mult_Buf[75].Weight_n = Wgt_1_761;
         Mult_Buf[76].Feature_n = FeatureBuf_762;
         Mult_Buf[76].Weight_n = Wgt_1_762;
         Mult_Buf[77].Feature_n = FeatureBuf_763;
         Mult_Buf[77].Weight_n = Wgt_1_763;
         Mult_Buf[78].Feature_n = FeatureBuf_764;
         Mult_Buf[78].Weight_n = Wgt_1_764;
         Mult_Buf[79].Feature_n = FeatureBuf_765;
         Mult_Buf[79].Weight_n = Wgt_1_765;
         Mult_Buf[80].Feature_n = FeatureBuf_766;
         Mult_Buf[80].Weight_n = Wgt_1_766;
         Mult_Buf[81].Feature_n = FeatureBuf_767;
         Mult_Buf[81].Weight_n = Wgt_1_767;
         Mult_Buf[82].Feature_n = FeatureBuf_768;
         Mult_Buf[82].Weight_n = Wgt_1_768;
         Mult_Buf[83].Feature_n = FeatureBuf_769;
         Mult_Buf[83].Weight_n = Wgt_1_769;
         Mult_Buf[84].Feature_n = FeatureBuf_770;
         Mult_Buf[84].Weight_n = Wgt_1_770;
         Mult_Buf[85].Feature_n = FeatureBuf_771;
         Mult_Buf[85].Weight_n = Wgt_1_771;
         Mult_Buf[86].Feature_n = FeatureBuf_772;
         Mult_Buf[86].Weight_n = Wgt_1_772;
         Mult_Buf[87].Feature_n = FeatureBuf_773;
         Mult_Buf[87].Weight_n = Wgt_1_773;
         Mult_Buf[88].Feature_n = FeatureBuf_774;
         Mult_Buf[88].Weight_n = Wgt_1_774;
         Mult_Buf[89].Feature_n = FeatureBuf_775;
         Mult_Buf[89].Weight_n = Wgt_1_775;
         Mult_Buf[90].Feature_n = FeatureBuf_776;
         Mult_Buf[90].Weight_n = Wgt_1_776;
         Mult_Buf[91].Feature_n = FeatureBuf_777;
         Mult_Buf[91].Weight_n = Wgt_1_777;
         Mult_Buf[92].Feature_n = FeatureBuf_778;
         Mult_Buf[92].Weight_n = Wgt_1_778;
         Mult_Buf[93].Feature_n = FeatureBuf_779;
         Mult_Buf[93].Weight_n = Wgt_1_779;
         Mult_Buf[94].Feature_n = FeatureBuf_780;
         Mult_Buf[94].Weight_n = Wgt_1_780;
         Mult_Buf[95].Feature_n = FeatureBuf_781;
         Mult_Buf[95].Weight_n = Wgt_1_781;
         Mult_Buf[96].Feature_n = FeatureBuf_782;
         Mult_Buf[96].Weight_n = Wgt_1_782;
         Mult_Buf[97].Feature_n = FeatureBuf_783;
         Mult_Buf[97].Weight_n = Wgt_1_783;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     end
    18:begin
     nxt_state = 19;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_0;
         Mult_Buf[0].Weight_n = Wgt_2_0;
         Mult_Buf[1].Feature_n = FeatureBuf_1;
         Mult_Buf[1].Weight_n = Wgt_2_1;
         Mult_Buf[2].Feature_n = FeatureBuf_2;
         Mult_Buf[2].Weight_n = Wgt_2_2;
         Mult_Buf[3].Feature_n = FeatureBuf_3;
         Mult_Buf[3].Weight_n = Wgt_2_3;
         Mult_Buf[4].Feature_n = FeatureBuf_4;
         Mult_Buf[4].Weight_n = Wgt_2_4;
         Mult_Buf[5].Feature_n = FeatureBuf_5;
         Mult_Buf[5].Weight_n = Wgt_2_5;
         Mult_Buf[6].Feature_n = FeatureBuf_6;
         Mult_Buf[6].Weight_n = Wgt_2_6;
         Mult_Buf[7].Feature_n = FeatureBuf_7;
         Mult_Buf[7].Weight_n = Wgt_2_7;
         Mult_Buf[8].Feature_n = FeatureBuf_8;
         Mult_Buf[8].Weight_n = Wgt_2_8;
         Mult_Buf[9].Feature_n = FeatureBuf_9;
         Mult_Buf[9].Weight_n = Wgt_2_9;
         Mult_Buf[10].Feature_n = FeatureBuf_10;
         Mult_Buf[10].Weight_n = Wgt_2_10;
         Mult_Buf[11].Feature_n = FeatureBuf_11;
         Mult_Buf[11].Weight_n = Wgt_2_11;
         Mult_Buf[12].Feature_n = FeatureBuf_12;
         Mult_Buf[12].Weight_n = Wgt_2_12;
         Mult_Buf[13].Feature_n = FeatureBuf_13;
         Mult_Buf[13].Weight_n = Wgt_2_13;
         Mult_Buf[14].Feature_n = FeatureBuf_14;
         Mult_Buf[14].Weight_n = Wgt_2_14;
         Mult_Buf[15].Feature_n = FeatureBuf_15;
         Mult_Buf[15].Weight_n = Wgt_2_15;
         Mult_Buf[16].Feature_n = FeatureBuf_16;
         Mult_Buf[16].Weight_n = Wgt_2_16;
         Mult_Buf[17].Feature_n = FeatureBuf_17;
         Mult_Buf[17].Weight_n = Wgt_2_17;
         Mult_Buf[18].Feature_n = FeatureBuf_18;
         Mult_Buf[18].Weight_n = Wgt_2_18;
         Mult_Buf[19].Feature_n = FeatureBuf_19;
         Mult_Buf[19].Weight_n = Wgt_2_19;
         Mult_Buf[20].Feature_n = FeatureBuf_20;
         Mult_Buf[20].Weight_n = Wgt_2_20;
         Mult_Buf[21].Feature_n = FeatureBuf_21;
         Mult_Buf[21].Weight_n = Wgt_2_21;
         Mult_Buf[22].Feature_n = FeatureBuf_22;
         Mult_Buf[22].Weight_n = Wgt_2_22;
         Mult_Buf[23].Feature_n = FeatureBuf_23;
         Mult_Buf[23].Weight_n = Wgt_2_23;
         Mult_Buf[24].Feature_n = FeatureBuf_24;
         Mult_Buf[24].Weight_n = Wgt_2_24;
         Mult_Buf[25].Feature_n = FeatureBuf_25;
         Mult_Buf[25].Weight_n = Wgt_2_25;
         Mult_Buf[26].Feature_n = FeatureBuf_26;
         Mult_Buf[26].Weight_n = Wgt_2_26;
         Mult_Buf[27].Feature_n = FeatureBuf_27;
         Mult_Buf[27].Weight_n = Wgt_2_27;
         Mult_Buf[28].Feature_n = FeatureBuf_28;
         Mult_Buf[28].Weight_n = Wgt_2_28;
         Mult_Buf[29].Feature_n = FeatureBuf_29;
         Mult_Buf[29].Weight_n = Wgt_2_29;
         Mult_Buf[30].Feature_n = FeatureBuf_30;
         Mult_Buf[30].Weight_n = Wgt_2_30;
         Mult_Buf[31].Feature_n = FeatureBuf_31;
         Mult_Buf[31].Weight_n = Wgt_2_31;
         Mult_Buf[32].Feature_n = FeatureBuf_32;
         Mult_Buf[32].Weight_n = Wgt_2_32;
         Mult_Buf[33].Feature_n = FeatureBuf_33;
         Mult_Buf[33].Weight_n = Wgt_2_33;
         Mult_Buf[34].Feature_n = FeatureBuf_34;
         Mult_Buf[34].Weight_n = Wgt_2_34;
         Mult_Buf[35].Feature_n = FeatureBuf_35;
         Mult_Buf[35].Weight_n = Wgt_2_35;
         Mult_Buf[36].Feature_n = FeatureBuf_36;
         Mult_Buf[36].Weight_n = Wgt_2_36;
         Mult_Buf[37].Feature_n = FeatureBuf_37;
         Mult_Buf[37].Weight_n = Wgt_2_37;
         Mult_Buf[38].Feature_n = FeatureBuf_38;
         Mult_Buf[38].Weight_n = Wgt_2_38;
         Mult_Buf[39].Feature_n = FeatureBuf_39;
         Mult_Buf[39].Weight_n = Wgt_2_39;
         Mult_Buf[40].Feature_n = FeatureBuf_40;
         Mult_Buf[40].Weight_n = Wgt_2_40;
         Mult_Buf[41].Feature_n = FeatureBuf_41;
         Mult_Buf[41].Weight_n = Wgt_2_41;
         Mult_Buf[42].Feature_n = FeatureBuf_42;
         Mult_Buf[42].Weight_n = Wgt_2_42;
         Mult_Buf[43].Feature_n = FeatureBuf_43;
         Mult_Buf[43].Weight_n = Wgt_2_43;
         Mult_Buf[44].Feature_n = FeatureBuf_44;
         Mult_Buf[44].Weight_n = Wgt_2_44;
         Mult_Buf[45].Feature_n = FeatureBuf_45;
         Mult_Buf[45].Weight_n = Wgt_2_45;
         Mult_Buf[46].Feature_n = FeatureBuf_46;
         Mult_Buf[46].Weight_n = Wgt_2_46;
         Mult_Buf[47].Feature_n = FeatureBuf_47;
         Mult_Buf[47].Weight_n = Wgt_2_47;
         Mult_Buf[48].Feature_n = FeatureBuf_48;
         Mult_Buf[48].Weight_n = Wgt_2_48;
         Mult_Buf[49].Feature_n = FeatureBuf_49;
         Mult_Buf[49].Weight_n = Wgt_2_49;
         Mult_Buf[50].Feature_n = FeatureBuf_50;
         Mult_Buf[50].Weight_n = Wgt_2_50;
         Mult_Buf[51].Feature_n = FeatureBuf_51;
         Mult_Buf[51].Weight_n = Wgt_2_51;
         Mult_Buf[52].Feature_n = FeatureBuf_52;
         Mult_Buf[52].Weight_n = Wgt_2_52;
         Mult_Buf[53].Feature_n = FeatureBuf_53;
         Mult_Buf[53].Weight_n = Wgt_2_53;
         Mult_Buf[54].Feature_n = FeatureBuf_54;
         Mult_Buf[54].Weight_n = Wgt_2_54;
         Mult_Buf[55].Feature_n = FeatureBuf_55;
         Mult_Buf[55].Weight_n = Wgt_2_55;
         Mult_Buf[56].Feature_n = FeatureBuf_56;
         Mult_Buf[56].Weight_n = Wgt_2_56;
         Mult_Buf[57].Feature_n = FeatureBuf_57;
         Mult_Buf[57].Weight_n = Wgt_2_57;
         Mult_Buf[58].Feature_n = FeatureBuf_58;
         Mult_Buf[58].Weight_n = Wgt_2_58;
         Mult_Buf[59].Feature_n = FeatureBuf_59;
         Mult_Buf[59].Weight_n = Wgt_2_59;
         Mult_Buf[60].Feature_n = FeatureBuf_60;
         Mult_Buf[60].Weight_n = Wgt_2_60;
         Mult_Buf[61].Feature_n = FeatureBuf_61;
         Mult_Buf[61].Weight_n = Wgt_2_61;
         Mult_Buf[62].Feature_n = FeatureBuf_62;
         Mult_Buf[62].Weight_n = Wgt_2_62;
         Mult_Buf[63].Feature_n = FeatureBuf_63;
         Mult_Buf[63].Weight_n = Wgt_2_63;
         Mult_Buf[64].Feature_n = FeatureBuf_64;
         Mult_Buf[64].Weight_n = Wgt_2_64;
         Mult_Buf[65].Feature_n = FeatureBuf_65;
         Mult_Buf[65].Weight_n = Wgt_2_65;
         Mult_Buf[66].Feature_n = FeatureBuf_66;
         Mult_Buf[66].Weight_n = Wgt_2_66;
         Mult_Buf[67].Feature_n = FeatureBuf_67;
         Mult_Buf[67].Weight_n = Wgt_2_67;
         Mult_Buf[68].Feature_n = FeatureBuf_68;
         Mult_Buf[68].Weight_n = Wgt_2_68;
         Mult_Buf[69].Feature_n = FeatureBuf_69;
         Mult_Buf[69].Weight_n = Wgt_2_69;
         Mult_Buf[70].Feature_n = FeatureBuf_70;
         Mult_Buf[70].Weight_n = Wgt_2_70;
         Mult_Buf[71].Feature_n = FeatureBuf_71;
         Mult_Buf[71].Weight_n = Wgt_2_71;
         Mult_Buf[72].Feature_n = FeatureBuf_72;
         Mult_Buf[72].Weight_n = Wgt_2_72;
         Mult_Buf[73].Feature_n = FeatureBuf_73;
         Mult_Buf[73].Weight_n = Wgt_2_73;
         Mult_Buf[74].Feature_n = FeatureBuf_74;
         Mult_Buf[74].Weight_n = Wgt_2_74;
         Mult_Buf[75].Feature_n = FeatureBuf_75;
         Mult_Buf[75].Weight_n = Wgt_2_75;
         Mult_Buf[76].Feature_n = FeatureBuf_76;
         Mult_Buf[76].Weight_n = Wgt_2_76;
         Mult_Buf[77].Feature_n = FeatureBuf_77;
         Mult_Buf[77].Weight_n = Wgt_2_77;
         Mult_Buf[78].Feature_n = FeatureBuf_78;
         Mult_Buf[78].Weight_n = Wgt_2_78;
         Mult_Buf[79].Feature_n = FeatureBuf_79;
         Mult_Buf[79].Weight_n = Wgt_2_79;
         Mult_Buf[80].Feature_n = FeatureBuf_80;
         Mult_Buf[80].Weight_n = Wgt_2_80;
         Mult_Buf[81].Feature_n = FeatureBuf_81;
         Mult_Buf[81].Weight_n = Wgt_2_81;
         Mult_Buf[82].Feature_n = FeatureBuf_82;
         Mult_Buf[82].Weight_n = Wgt_2_82;
         Mult_Buf[83].Feature_n = FeatureBuf_83;
         Mult_Buf[83].Weight_n = Wgt_2_83;
         Mult_Buf[84].Feature_n = FeatureBuf_84;
         Mult_Buf[84].Weight_n = Wgt_2_84;
         Mult_Buf[85].Feature_n = FeatureBuf_85;
         Mult_Buf[85].Weight_n = Wgt_2_85;
         Mult_Buf[86].Feature_n = FeatureBuf_86;
         Mult_Buf[86].Weight_n = Wgt_2_86;
         Mult_Buf[87].Feature_n = FeatureBuf_87;
         Mult_Buf[87].Weight_n = Wgt_2_87;
         Mult_Buf[88].Feature_n = FeatureBuf_88;
         Mult_Buf[88].Weight_n = Wgt_2_88;
         Mult_Buf[89].Feature_n = FeatureBuf_89;
         Mult_Buf[89].Weight_n = Wgt_2_89;
         Mult_Buf[90].Feature_n = FeatureBuf_90;
         Mult_Buf[90].Weight_n = Wgt_2_90;
         Mult_Buf[91].Feature_n = FeatureBuf_91;
         Mult_Buf[91].Weight_n = Wgt_2_91;
         Mult_Buf[92].Feature_n = FeatureBuf_92;
         Mult_Buf[92].Weight_n = Wgt_2_92;
         Mult_Buf[93].Feature_n = FeatureBuf_93;
         Mult_Buf[93].Weight_n = Wgt_2_93;
         Mult_Buf[94].Feature_n = FeatureBuf_94;
         Mult_Buf[94].Weight_n = Wgt_2_94;
         Mult_Buf[95].Feature_n = FeatureBuf_95;
         Mult_Buf[95].Weight_n = Wgt_2_95;
         Mult_Buf[96].Feature_n = FeatureBuf_96;
         Mult_Buf[96].Weight_n = Wgt_2_96;
         Mult_Buf[97].Feature_n = FeatureBuf_97;
         Mult_Buf[97].Weight_n = Wgt_2_97;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     end
    19:begin
     nxt_state = 20;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_98;
         Mult_Buf[0].Weight_n = Wgt_2_98;
         Mult_Buf[1].Feature_n = FeatureBuf_99;
         Mult_Buf[1].Weight_n = Wgt_2_99;
         Mult_Buf[2].Feature_n = FeatureBuf_100;
         Mult_Buf[2].Weight_n = Wgt_2_100;
         Mult_Buf[3].Feature_n = FeatureBuf_101;
         Mult_Buf[3].Weight_n = Wgt_2_101;
         Mult_Buf[4].Feature_n = FeatureBuf_102;
         Mult_Buf[4].Weight_n = Wgt_2_102;
         Mult_Buf[5].Feature_n = FeatureBuf_103;
         Mult_Buf[5].Weight_n = Wgt_2_103;
         Mult_Buf[6].Feature_n = FeatureBuf_104;
         Mult_Buf[6].Weight_n = Wgt_2_104;
         Mult_Buf[7].Feature_n = FeatureBuf_105;
         Mult_Buf[7].Weight_n = Wgt_2_105;
         Mult_Buf[8].Feature_n = FeatureBuf_106;
         Mult_Buf[8].Weight_n = Wgt_2_106;
         Mult_Buf[9].Feature_n = FeatureBuf_107;
         Mult_Buf[9].Weight_n = Wgt_2_107;
         Mult_Buf[10].Feature_n = FeatureBuf_108;
         Mult_Buf[10].Weight_n = Wgt_2_108;
         Mult_Buf[11].Feature_n = FeatureBuf_109;
         Mult_Buf[11].Weight_n = Wgt_2_109;
         Mult_Buf[12].Feature_n = FeatureBuf_110;
         Mult_Buf[12].Weight_n = Wgt_2_110;
         Mult_Buf[13].Feature_n = FeatureBuf_111;
         Mult_Buf[13].Weight_n = Wgt_2_111;
         Mult_Buf[14].Feature_n = FeatureBuf_112;
         Mult_Buf[14].Weight_n = Wgt_2_112;
         Mult_Buf[15].Feature_n = FeatureBuf_113;
         Mult_Buf[15].Weight_n = Wgt_2_113;
         Mult_Buf[16].Feature_n = FeatureBuf_114;
         Mult_Buf[16].Weight_n = Wgt_2_114;
         Mult_Buf[17].Feature_n = FeatureBuf_115;
         Mult_Buf[17].Weight_n = Wgt_2_115;
         Mult_Buf[18].Feature_n = FeatureBuf_116;
         Mult_Buf[18].Weight_n = Wgt_2_116;
         Mult_Buf[19].Feature_n = FeatureBuf_117;
         Mult_Buf[19].Weight_n = Wgt_2_117;
         Mult_Buf[20].Feature_n = FeatureBuf_118;
         Mult_Buf[20].Weight_n = Wgt_2_118;
         Mult_Buf[21].Feature_n = FeatureBuf_119;
         Mult_Buf[21].Weight_n = Wgt_2_119;
         Mult_Buf[22].Feature_n = FeatureBuf_120;
         Mult_Buf[22].Weight_n = Wgt_2_120;
         Mult_Buf[23].Feature_n = FeatureBuf_121;
         Mult_Buf[23].Weight_n = Wgt_2_121;
         Mult_Buf[24].Feature_n = FeatureBuf_122;
         Mult_Buf[24].Weight_n = Wgt_2_122;
         Mult_Buf[25].Feature_n = FeatureBuf_123;
         Mult_Buf[25].Weight_n = Wgt_2_123;
         Mult_Buf[26].Feature_n = FeatureBuf_124;
         Mult_Buf[26].Weight_n = Wgt_2_124;
         Mult_Buf[27].Feature_n = FeatureBuf_125;
         Mult_Buf[27].Weight_n = Wgt_2_125;
         Mult_Buf[28].Feature_n = FeatureBuf_126;
         Mult_Buf[28].Weight_n = Wgt_2_126;
         Mult_Buf[29].Feature_n = FeatureBuf_127;
         Mult_Buf[29].Weight_n = Wgt_2_127;
         Mult_Buf[30].Feature_n = FeatureBuf_128;
         Mult_Buf[30].Weight_n = Wgt_2_128;
         Mult_Buf[31].Feature_n = FeatureBuf_129;
         Mult_Buf[31].Weight_n = Wgt_2_129;
         Mult_Buf[32].Feature_n = FeatureBuf_130;
         Mult_Buf[32].Weight_n = Wgt_2_130;
         Mult_Buf[33].Feature_n = FeatureBuf_131;
         Mult_Buf[33].Weight_n = Wgt_2_131;
         Mult_Buf[34].Feature_n = FeatureBuf_132;
         Mult_Buf[34].Weight_n = Wgt_2_132;
         Mult_Buf[35].Feature_n = FeatureBuf_133;
         Mult_Buf[35].Weight_n = Wgt_2_133;
         Mult_Buf[36].Feature_n = FeatureBuf_134;
         Mult_Buf[36].Weight_n = Wgt_2_134;
         Mult_Buf[37].Feature_n = FeatureBuf_135;
         Mult_Buf[37].Weight_n = Wgt_2_135;
         Mult_Buf[38].Feature_n = FeatureBuf_136;
         Mult_Buf[38].Weight_n = Wgt_2_136;
         Mult_Buf[39].Feature_n = FeatureBuf_137;
         Mult_Buf[39].Weight_n = Wgt_2_137;
         Mult_Buf[40].Feature_n = FeatureBuf_138;
         Mult_Buf[40].Weight_n = Wgt_2_138;
         Mult_Buf[41].Feature_n = FeatureBuf_139;
         Mult_Buf[41].Weight_n = Wgt_2_139;
         Mult_Buf[42].Feature_n = FeatureBuf_140;
         Mult_Buf[42].Weight_n = Wgt_2_140;
         Mult_Buf[43].Feature_n = FeatureBuf_141;
         Mult_Buf[43].Weight_n = Wgt_2_141;
         Mult_Buf[44].Feature_n = FeatureBuf_142;
         Mult_Buf[44].Weight_n = Wgt_2_142;
         Mult_Buf[45].Feature_n = FeatureBuf_143;
         Mult_Buf[45].Weight_n = Wgt_2_143;
         Mult_Buf[46].Feature_n = FeatureBuf_144;
         Mult_Buf[46].Weight_n = Wgt_2_144;
         Mult_Buf[47].Feature_n = FeatureBuf_145;
         Mult_Buf[47].Weight_n = Wgt_2_145;
         Mult_Buf[48].Feature_n = FeatureBuf_146;
         Mult_Buf[48].Weight_n = Wgt_2_146;
         Mult_Buf[49].Feature_n = FeatureBuf_147;
         Mult_Buf[49].Weight_n = Wgt_2_147;
         Mult_Buf[50].Feature_n = FeatureBuf_148;
         Mult_Buf[50].Weight_n = Wgt_2_148;
         Mult_Buf[51].Feature_n = FeatureBuf_149;
         Mult_Buf[51].Weight_n = Wgt_2_149;
         Mult_Buf[52].Feature_n = FeatureBuf_150;
         Mult_Buf[52].Weight_n = Wgt_2_150;
         Mult_Buf[53].Feature_n = FeatureBuf_151;
         Mult_Buf[53].Weight_n = Wgt_2_151;
         Mult_Buf[54].Feature_n = FeatureBuf_152;
         Mult_Buf[54].Weight_n = Wgt_2_152;
         Mult_Buf[55].Feature_n = FeatureBuf_153;
         Mult_Buf[55].Weight_n = Wgt_2_153;
         Mult_Buf[56].Feature_n = FeatureBuf_154;
         Mult_Buf[56].Weight_n = Wgt_2_154;
         Mult_Buf[57].Feature_n = FeatureBuf_155;
         Mult_Buf[57].Weight_n = Wgt_2_155;
         Mult_Buf[58].Feature_n = FeatureBuf_156;
         Mult_Buf[58].Weight_n = Wgt_2_156;
         Mult_Buf[59].Feature_n = FeatureBuf_157;
         Mult_Buf[59].Weight_n = Wgt_2_157;
         Mult_Buf[60].Feature_n = FeatureBuf_158;
         Mult_Buf[60].Weight_n = Wgt_2_158;
         Mult_Buf[61].Feature_n = FeatureBuf_159;
         Mult_Buf[61].Weight_n = Wgt_2_159;
         Mult_Buf[62].Feature_n = FeatureBuf_160;
         Mult_Buf[62].Weight_n = Wgt_2_160;
         Mult_Buf[63].Feature_n = FeatureBuf_161;
         Mult_Buf[63].Weight_n = Wgt_2_161;
         Mult_Buf[64].Feature_n = FeatureBuf_162;
         Mult_Buf[64].Weight_n = Wgt_2_162;
         Mult_Buf[65].Feature_n = FeatureBuf_163;
         Mult_Buf[65].Weight_n = Wgt_2_163;
         Mult_Buf[66].Feature_n = FeatureBuf_164;
         Mult_Buf[66].Weight_n = Wgt_2_164;
         Mult_Buf[67].Feature_n = FeatureBuf_165;
         Mult_Buf[67].Weight_n = Wgt_2_165;
         Mult_Buf[68].Feature_n = FeatureBuf_166;
         Mult_Buf[68].Weight_n = Wgt_2_166;
         Mult_Buf[69].Feature_n = FeatureBuf_167;
         Mult_Buf[69].Weight_n = Wgt_2_167;
         Mult_Buf[70].Feature_n = FeatureBuf_168;
         Mult_Buf[70].Weight_n = Wgt_2_168;
         Mult_Buf[71].Feature_n = FeatureBuf_169;
         Mult_Buf[71].Weight_n = Wgt_2_169;
         Mult_Buf[72].Feature_n = FeatureBuf_170;
         Mult_Buf[72].Weight_n = Wgt_2_170;
         Mult_Buf[73].Feature_n = FeatureBuf_171;
         Mult_Buf[73].Weight_n = Wgt_2_171;
         Mult_Buf[74].Feature_n = FeatureBuf_172;
         Mult_Buf[74].Weight_n = Wgt_2_172;
         Mult_Buf[75].Feature_n = FeatureBuf_173;
         Mult_Buf[75].Weight_n = Wgt_2_173;
         Mult_Buf[76].Feature_n = FeatureBuf_174;
         Mult_Buf[76].Weight_n = Wgt_2_174;
         Mult_Buf[77].Feature_n = FeatureBuf_175;
         Mult_Buf[77].Weight_n = Wgt_2_175;
         Mult_Buf[78].Feature_n = FeatureBuf_176;
         Mult_Buf[78].Weight_n = Wgt_2_176;
         Mult_Buf[79].Feature_n = FeatureBuf_177;
         Mult_Buf[79].Weight_n = Wgt_2_177;
         Mult_Buf[80].Feature_n = FeatureBuf_178;
         Mult_Buf[80].Weight_n = Wgt_2_178;
         Mult_Buf[81].Feature_n = FeatureBuf_179;
         Mult_Buf[81].Weight_n = Wgt_2_179;
         Mult_Buf[82].Feature_n = FeatureBuf_180;
         Mult_Buf[82].Weight_n = Wgt_2_180;
         Mult_Buf[83].Feature_n = FeatureBuf_181;
         Mult_Buf[83].Weight_n = Wgt_2_181;
         Mult_Buf[84].Feature_n = FeatureBuf_182;
         Mult_Buf[84].Weight_n = Wgt_2_182;
         Mult_Buf[85].Feature_n = FeatureBuf_183;
         Mult_Buf[85].Weight_n = Wgt_2_183;
         Mult_Buf[86].Feature_n = FeatureBuf_184;
         Mult_Buf[86].Weight_n = Wgt_2_184;
         Mult_Buf[87].Feature_n = FeatureBuf_185;
         Mult_Buf[87].Weight_n = Wgt_2_185;
         Mult_Buf[88].Feature_n = FeatureBuf_186;
         Mult_Buf[88].Weight_n = Wgt_2_186;
         Mult_Buf[89].Feature_n = FeatureBuf_187;
         Mult_Buf[89].Weight_n = Wgt_2_187;
         Mult_Buf[90].Feature_n = FeatureBuf_188;
         Mult_Buf[90].Weight_n = Wgt_2_188;
         Mult_Buf[91].Feature_n = FeatureBuf_189;
         Mult_Buf[91].Weight_n = Wgt_2_189;
         Mult_Buf[92].Feature_n = FeatureBuf_190;
         Mult_Buf[92].Weight_n = Wgt_2_190;
         Mult_Buf[93].Feature_n = FeatureBuf_191;
         Mult_Buf[93].Weight_n = Wgt_2_191;
         Mult_Buf[94].Feature_n = FeatureBuf_192;
         Mult_Buf[94].Weight_n = Wgt_2_192;
         Mult_Buf[95].Feature_n = FeatureBuf_193;
         Mult_Buf[95].Weight_n = Wgt_2_193;
         Mult_Buf[96].Feature_n = FeatureBuf_194;
         Mult_Buf[96].Weight_n = Wgt_2_194;
         Mult_Buf[97].Feature_n = FeatureBuf_195;
         Mult_Buf[97].Weight_n = Wgt_2_195;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     end
    20:begin
     nxt_state = 21;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_196;
         Mult_Buf[0].Weight_n = Wgt_2_196;
         Mult_Buf[1].Feature_n = FeatureBuf_197;
         Mult_Buf[1].Weight_n = Wgt_2_197;
         Mult_Buf[2].Feature_n = FeatureBuf_198;
         Mult_Buf[2].Weight_n = Wgt_2_198;
         Mult_Buf[3].Feature_n = FeatureBuf_199;
         Mult_Buf[3].Weight_n = Wgt_2_199;
         Mult_Buf[4].Feature_n = FeatureBuf_200;
         Mult_Buf[4].Weight_n = Wgt_2_200;
         Mult_Buf[5].Feature_n = FeatureBuf_201;
         Mult_Buf[5].Weight_n = Wgt_2_201;
         Mult_Buf[6].Feature_n = FeatureBuf_202;
         Mult_Buf[6].Weight_n = Wgt_2_202;
         Mult_Buf[7].Feature_n = FeatureBuf_203;
         Mult_Buf[7].Weight_n = Wgt_2_203;
         Mult_Buf[8].Feature_n = FeatureBuf_204;
         Mult_Buf[8].Weight_n = Wgt_2_204;
         Mult_Buf[9].Feature_n = FeatureBuf_205;
         Mult_Buf[9].Weight_n = Wgt_2_205;
         Mult_Buf[10].Feature_n = FeatureBuf_206;
         Mult_Buf[10].Weight_n = Wgt_2_206;
         Mult_Buf[11].Feature_n = FeatureBuf_207;
         Mult_Buf[11].Weight_n = Wgt_2_207;
         Mult_Buf[12].Feature_n = FeatureBuf_208;
         Mult_Buf[12].Weight_n = Wgt_2_208;
         Mult_Buf[13].Feature_n = FeatureBuf_209;
         Mult_Buf[13].Weight_n = Wgt_2_209;
         Mult_Buf[14].Feature_n = FeatureBuf_210;
         Mult_Buf[14].Weight_n = Wgt_2_210;
         Mult_Buf[15].Feature_n = FeatureBuf_211;
         Mult_Buf[15].Weight_n = Wgt_2_211;
         Mult_Buf[16].Feature_n = FeatureBuf_212;
         Mult_Buf[16].Weight_n = Wgt_2_212;
         Mult_Buf[17].Feature_n = FeatureBuf_213;
         Mult_Buf[17].Weight_n = Wgt_2_213;
         Mult_Buf[18].Feature_n = FeatureBuf_214;
         Mult_Buf[18].Weight_n = Wgt_2_214;
         Mult_Buf[19].Feature_n = FeatureBuf_215;
         Mult_Buf[19].Weight_n = Wgt_2_215;
         Mult_Buf[20].Feature_n = FeatureBuf_216;
         Mult_Buf[20].Weight_n = Wgt_2_216;
         Mult_Buf[21].Feature_n = FeatureBuf_217;
         Mult_Buf[21].Weight_n = Wgt_2_217;
         Mult_Buf[22].Feature_n = FeatureBuf_218;
         Mult_Buf[22].Weight_n = Wgt_2_218;
         Mult_Buf[23].Feature_n = FeatureBuf_219;
         Mult_Buf[23].Weight_n = Wgt_2_219;
         Mult_Buf[24].Feature_n = FeatureBuf_220;
         Mult_Buf[24].Weight_n = Wgt_2_220;
         Mult_Buf[25].Feature_n = FeatureBuf_221;
         Mult_Buf[25].Weight_n = Wgt_2_221;
         Mult_Buf[26].Feature_n = FeatureBuf_222;
         Mult_Buf[26].Weight_n = Wgt_2_222;
         Mult_Buf[27].Feature_n = FeatureBuf_223;
         Mult_Buf[27].Weight_n = Wgt_2_223;
         Mult_Buf[28].Feature_n = FeatureBuf_224;
         Mult_Buf[28].Weight_n = Wgt_2_224;
         Mult_Buf[29].Feature_n = FeatureBuf_225;
         Mult_Buf[29].Weight_n = Wgt_2_225;
         Mult_Buf[30].Feature_n = FeatureBuf_226;
         Mult_Buf[30].Weight_n = Wgt_2_226;
         Mult_Buf[31].Feature_n = FeatureBuf_227;
         Mult_Buf[31].Weight_n = Wgt_2_227;
         Mult_Buf[32].Feature_n = FeatureBuf_228;
         Mult_Buf[32].Weight_n = Wgt_2_228;
         Mult_Buf[33].Feature_n = FeatureBuf_229;
         Mult_Buf[33].Weight_n = Wgt_2_229;
         Mult_Buf[34].Feature_n = FeatureBuf_230;
         Mult_Buf[34].Weight_n = Wgt_2_230;
         Mult_Buf[35].Feature_n = FeatureBuf_231;
         Mult_Buf[35].Weight_n = Wgt_2_231;
         Mult_Buf[36].Feature_n = FeatureBuf_232;
         Mult_Buf[36].Weight_n = Wgt_2_232;
         Mult_Buf[37].Feature_n = FeatureBuf_233;
         Mult_Buf[37].Weight_n = Wgt_2_233;
         Mult_Buf[38].Feature_n = FeatureBuf_234;
         Mult_Buf[38].Weight_n = Wgt_2_234;
         Mult_Buf[39].Feature_n = FeatureBuf_235;
         Mult_Buf[39].Weight_n = Wgt_2_235;
         Mult_Buf[40].Feature_n = FeatureBuf_236;
         Mult_Buf[40].Weight_n = Wgt_2_236;
         Mult_Buf[41].Feature_n = FeatureBuf_237;
         Mult_Buf[41].Weight_n = Wgt_2_237;
         Mult_Buf[42].Feature_n = FeatureBuf_238;
         Mult_Buf[42].Weight_n = Wgt_2_238;
         Mult_Buf[43].Feature_n = FeatureBuf_239;
         Mult_Buf[43].Weight_n = Wgt_2_239;
         Mult_Buf[44].Feature_n = FeatureBuf_240;
         Mult_Buf[44].Weight_n = Wgt_2_240;
         Mult_Buf[45].Feature_n = FeatureBuf_241;
         Mult_Buf[45].Weight_n = Wgt_2_241;
         Mult_Buf[46].Feature_n = FeatureBuf_242;
         Mult_Buf[46].Weight_n = Wgt_2_242;
         Mult_Buf[47].Feature_n = FeatureBuf_243;
         Mult_Buf[47].Weight_n = Wgt_2_243;
         Mult_Buf[48].Feature_n = FeatureBuf_244;
         Mult_Buf[48].Weight_n = Wgt_2_244;
         Mult_Buf[49].Feature_n = FeatureBuf_245;
         Mult_Buf[49].Weight_n = Wgt_2_245;
         Mult_Buf[50].Feature_n = FeatureBuf_246;
         Mult_Buf[50].Weight_n = Wgt_2_246;
         Mult_Buf[51].Feature_n = FeatureBuf_247;
         Mult_Buf[51].Weight_n = Wgt_2_247;
         Mult_Buf[52].Feature_n = FeatureBuf_248;
         Mult_Buf[52].Weight_n = Wgt_2_248;
         Mult_Buf[53].Feature_n = FeatureBuf_249;
         Mult_Buf[53].Weight_n = Wgt_2_249;
         Mult_Buf[54].Feature_n = FeatureBuf_250;
         Mult_Buf[54].Weight_n = Wgt_2_250;
         Mult_Buf[55].Feature_n = FeatureBuf_251;
         Mult_Buf[55].Weight_n = Wgt_2_251;
         Mult_Buf[56].Feature_n = FeatureBuf_252;
         Mult_Buf[56].Weight_n = Wgt_2_252;
         Mult_Buf[57].Feature_n = FeatureBuf_253;
         Mult_Buf[57].Weight_n = Wgt_2_253;
         Mult_Buf[58].Feature_n = FeatureBuf_254;
         Mult_Buf[58].Weight_n = Wgt_2_254;
         Mult_Buf[59].Feature_n = FeatureBuf_255;
         Mult_Buf[59].Weight_n = Wgt_2_255;
         Mult_Buf[60].Feature_n = FeatureBuf_256;
         Mult_Buf[60].Weight_n = Wgt_2_256;
         Mult_Buf[61].Feature_n = FeatureBuf_257;
         Mult_Buf[61].Weight_n = Wgt_2_257;
         Mult_Buf[62].Feature_n = FeatureBuf_258;
         Mult_Buf[62].Weight_n = Wgt_2_258;
         Mult_Buf[63].Feature_n = FeatureBuf_259;
         Mult_Buf[63].Weight_n = Wgt_2_259;
         Mult_Buf[64].Feature_n = FeatureBuf_260;
         Mult_Buf[64].Weight_n = Wgt_2_260;
         Mult_Buf[65].Feature_n = FeatureBuf_261;
         Mult_Buf[65].Weight_n = Wgt_2_261;
         Mult_Buf[66].Feature_n = FeatureBuf_262;
         Mult_Buf[66].Weight_n = Wgt_2_262;
         Mult_Buf[67].Feature_n = FeatureBuf_263;
         Mult_Buf[67].Weight_n = Wgt_2_263;
         Mult_Buf[68].Feature_n = FeatureBuf_264;
         Mult_Buf[68].Weight_n = Wgt_2_264;
         Mult_Buf[69].Feature_n = FeatureBuf_265;
         Mult_Buf[69].Weight_n = Wgt_2_265;
         Mult_Buf[70].Feature_n = FeatureBuf_266;
         Mult_Buf[70].Weight_n = Wgt_2_266;
         Mult_Buf[71].Feature_n = FeatureBuf_267;
         Mult_Buf[71].Weight_n = Wgt_2_267;
         Mult_Buf[72].Feature_n = FeatureBuf_268;
         Mult_Buf[72].Weight_n = Wgt_2_268;
         Mult_Buf[73].Feature_n = FeatureBuf_269;
         Mult_Buf[73].Weight_n = Wgt_2_269;
         Mult_Buf[74].Feature_n = FeatureBuf_270;
         Mult_Buf[74].Weight_n = Wgt_2_270;
         Mult_Buf[75].Feature_n = FeatureBuf_271;
         Mult_Buf[75].Weight_n = Wgt_2_271;
         Mult_Buf[76].Feature_n = FeatureBuf_272;
         Mult_Buf[76].Weight_n = Wgt_2_272;
         Mult_Buf[77].Feature_n = FeatureBuf_273;
         Mult_Buf[77].Weight_n = Wgt_2_273;
         Mult_Buf[78].Feature_n = FeatureBuf_274;
         Mult_Buf[78].Weight_n = Wgt_2_274;
         Mult_Buf[79].Feature_n = FeatureBuf_275;
         Mult_Buf[79].Weight_n = Wgt_2_275;
         Mult_Buf[80].Feature_n = FeatureBuf_276;
         Mult_Buf[80].Weight_n = Wgt_2_276;
         Mult_Buf[81].Feature_n = FeatureBuf_277;
         Mult_Buf[81].Weight_n = Wgt_2_277;
         Mult_Buf[82].Feature_n = FeatureBuf_278;
         Mult_Buf[82].Weight_n = Wgt_2_278;
         Mult_Buf[83].Feature_n = FeatureBuf_279;
         Mult_Buf[83].Weight_n = Wgt_2_279;
         Mult_Buf[84].Feature_n = FeatureBuf_280;
         Mult_Buf[84].Weight_n = Wgt_2_280;
         Mult_Buf[85].Feature_n = FeatureBuf_281;
         Mult_Buf[85].Weight_n = Wgt_2_281;
         Mult_Buf[86].Feature_n = FeatureBuf_282;
         Mult_Buf[86].Weight_n = Wgt_2_282;
         Mult_Buf[87].Feature_n = FeatureBuf_283;
         Mult_Buf[87].Weight_n = Wgt_2_283;
         Mult_Buf[88].Feature_n = FeatureBuf_284;
         Mult_Buf[88].Weight_n = Wgt_2_284;
         Mult_Buf[89].Feature_n = FeatureBuf_285;
         Mult_Buf[89].Weight_n = Wgt_2_285;
         Mult_Buf[90].Feature_n = FeatureBuf_286;
         Mult_Buf[90].Weight_n = Wgt_2_286;
         Mult_Buf[91].Feature_n = FeatureBuf_287;
         Mult_Buf[91].Weight_n = Wgt_2_287;
         Mult_Buf[92].Feature_n = FeatureBuf_288;
         Mult_Buf[92].Weight_n = Wgt_2_288;
         Mult_Buf[93].Feature_n = FeatureBuf_289;
         Mult_Buf[93].Weight_n = Wgt_2_289;
         Mult_Buf[94].Feature_n = FeatureBuf_290;
         Mult_Buf[94].Weight_n = Wgt_2_290;
         Mult_Buf[95].Feature_n = FeatureBuf_291;
         Mult_Buf[95].Weight_n = Wgt_2_291;
         Mult_Buf[96].Feature_n = FeatureBuf_292;
         Mult_Buf[96].Weight_n = Wgt_2_292;
         Mult_Buf[97].Feature_n = FeatureBuf_293;
         Mult_Buf[97].Weight_n = Wgt_2_293;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     end
    21:begin
     nxt_state = 22;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_294;
         Mult_Buf[0].Weight_n = Wgt_2_294;
         Mult_Buf[1].Feature_n = FeatureBuf_295;
         Mult_Buf[1].Weight_n = Wgt_2_295;
         Mult_Buf[2].Feature_n = FeatureBuf_296;
         Mult_Buf[2].Weight_n = Wgt_2_296;
         Mult_Buf[3].Feature_n = FeatureBuf_297;
         Mult_Buf[3].Weight_n = Wgt_2_297;
         Mult_Buf[4].Feature_n = FeatureBuf_298;
         Mult_Buf[4].Weight_n = Wgt_2_298;
         Mult_Buf[5].Feature_n = FeatureBuf_299;
         Mult_Buf[5].Weight_n = Wgt_2_299;
         Mult_Buf[6].Feature_n = FeatureBuf_300;
         Mult_Buf[6].Weight_n = Wgt_2_300;
         Mult_Buf[7].Feature_n = FeatureBuf_301;
         Mult_Buf[7].Weight_n = Wgt_2_301;
         Mult_Buf[8].Feature_n = FeatureBuf_302;
         Mult_Buf[8].Weight_n = Wgt_2_302;
         Mult_Buf[9].Feature_n = FeatureBuf_303;
         Mult_Buf[9].Weight_n = Wgt_2_303;
         Mult_Buf[10].Feature_n = FeatureBuf_304;
         Mult_Buf[10].Weight_n = Wgt_2_304;
         Mult_Buf[11].Feature_n = FeatureBuf_305;
         Mult_Buf[11].Weight_n = Wgt_2_305;
         Mult_Buf[12].Feature_n = FeatureBuf_306;
         Mult_Buf[12].Weight_n = Wgt_2_306;
         Mult_Buf[13].Feature_n = FeatureBuf_307;
         Mult_Buf[13].Weight_n = Wgt_2_307;
         Mult_Buf[14].Feature_n = FeatureBuf_308;
         Mult_Buf[14].Weight_n = Wgt_2_308;
         Mult_Buf[15].Feature_n = FeatureBuf_309;
         Mult_Buf[15].Weight_n = Wgt_2_309;
         Mult_Buf[16].Feature_n = FeatureBuf_310;
         Mult_Buf[16].Weight_n = Wgt_2_310;
         Mult_Buf[17].Feature_n = FeatureBuf_311;
         Mult_Buf[17].Weight_n = Wgt_2_311;
         Mult_Buf[18].Feature_n = FeatureBuf_312;
         Mult_Buf[18].Weight_n = Wgt_2_312;
         Mult_Buf[19].Feature_n = FeatureBuf_313;
         Mult_Buf[19].Weight_n = Wgt_2_313;
         Mult_Buf[20].Feature_n = FeatureBuf_314;
         Mult_Buf[20].Weight_n = Wgt_2_314;
         Mult_Buf[21].Feature_n = FeatureBuf_315;
         Mult_Buf[21].Weight_n = Wgt_2_315;
         Mult_Buf[22].Feature_n = FeatureBuf_316;
         Mult_Buf[22].Weight_n = Wgt_2_316;
         Mult_Buf[23].Feature_n = FeatureBuf_317;
         Mult_Buf[23].Weight_n = Wgt_2_317;
         Mult_Buf[24].Feature_n = FeatureBuf_318;
         Mult_Buf[24].Weight_n = Wgt_2_318;
         Mult_Buf[25].Feature_n = FeatureBuf_319;
         Mult_Buf[25].Weight_n = Wgt_2_319;
         Mult_Buf[26].Feature_n = FeatureBuf_320;
         Mult_Buf[26].Weight_n = Wgt_2_320;
         Mult_Buf[27].Feature_n = FeatureBuf_321;
         Mult_Buf[27].Weight_n = Wgt_2_321;
         Mult_Buf[28].Feature_n = FeatureBuf_322;
         Mult_Buf[28].Weight_n = Wgt_2_322;
         Mult_Buf[29].Feature_n = FeatureBuf_323;
         Mult_Buf[29].Weight_n = Wgt_2_323;
         Mult_Buf[30].Feature_n = FeatureBuf_324;
         Mult_Buf[30].Weight_n = Wgt_2_324;
         Mult_Buf[31].Feature_n = FeatureBuf_325;
         Mult_Buf[31].Weight_n = Wgt_2_325;
         Mult_Buf[32].Feature_n = FeatureBuf_326;
         Mult_Buf[32].Weight_n = Wgt_2_326;
         Mult_Buf[33].Feature_n = FeatureBuf_327;
         Mult_Buf[33].Weight_n = Wgt_2_327;
         Mult_Buf[34].Feature_n = FeatureBuf_328;
         Mult_Buf[34].Weight_n = Wgt_2_328;
         Mult_Buf[35].Feature_n = FeatureBuf_329;
         Mult_Buf[35].Weight_n = Wgt_2_329;
         Mult_Buf[36].Feature_n = FeatureBuf_330;
         Mult_Buf[36].Weight_n = Wgt_2_330;
         Mult_Buf[37].Feature_n = FeatureBuf_331;
         Mult_Buf[37].Weight_n = Wgt_2_331;
         Mult_Buf[38].Feature_n = FeatureBuf_332;
         Mult_Buf[38].Weight_n = Wgt_2_332;
         Mult_Buf[39].Feature_n = FeatureBuf_333;
         Mult_Buf[39].Weight_n = Wgt_2_333;
         Mult_Buf[40].Feature_n = FeatureBuf_334;
         Mult_Buf[40].Weight_n = Wgt_2_334;
         Mult_Buf[41].Feature_n = FeatureBuf_335;
         Mult_Buf[41].Weight_n = Wgt_2_335;
         Mult_Buf[42].Feature_n = FeatureBuf_336;
         Mult_Buf[42].Weight_n = Wgt_2_336;
         Mult_Buf[43].Feature_n = FeatureBuf_337;
         Mult_Buf[43].Weight_n = Wgt_2_337;
         Mult_Buf[44].Feature_n = FeatureBuf_338;
         Mult_Buf[44].Weight_n = Wgt_2_338;
         Mult_Buf[45].Feature_n = FeatureBuf_339;
         Mult_Buf[45].Weight_n = Wgt_2_339;
         Mult_Buf[46].Feature_n = FeatureBuf_340;
         Mult_Buf[46].Weight_n = Wgt_2_340;
         Mult_Buf[47].Feature_n = FeatureBuf_341;
         Mult_Buf[47].Weight_n = Wgt_2_341;
         Mult_Buf[48].Feature_n = FeatureBuf_342;
         Mult_Buf[48].Weight_n = Wgt_2_342;
         Mult_Buf[49].Feature_n = FeatureBuf_343;
         Mult_Buf[49].Weight_n = Wgt_2_343;
         Mult_Buf[50].Feature_n = FeatureBuf_344;
         Mult_Buf[50].Weight_n = Wgt_2_344;
         Mult_Buf[51].Feature_n = FeatureBuf_345;
         Mult_Buf[51].Weight_n = Wgt_2_345;
         Mult_Buf[52].Feature_n = FeatureBuf_346;
         Mult_Buf[52].Weight_n = Wgt_2_346;
         Mult_Buf[53].Feature_n = FeatureBuf_347;
         Mult_Buf[53].Weight_n = Wgt_2_347;
         Mult_Buf[54].Feature_n = FeatureBuf_348;
         Mult_Buf[54].Weight_n = Wgt_2_348;
         Mult_Buf[55].Feature_n = FeatureBuf_349;
         Mult_Buf[55].Weight_n = Wgt_2_349;
         Mult_Buf[56].Feature_n = FeatureBuf_350;
         Mult_Buf[56].Weight_n = Wgt_2_350;
         Mult_Buf[57].Feature_n = FeatureBuf_351;
         Mult_Buf[57].Weight_n = Wgt_2_351;
         Mult_Buf[58].Feature_n = FeatureBuf_352;
         Mult_Buf[58].Weight_n = Wgt_2_352;
         Mult_Buf[59].Feature_n = FeatureBuf_353;
         Mult_Buf[59].Weight_n = Wgt_2_353;
         Mult_Buf[60].Feature_n = FeatureBuf_354;
         Mult_Buf[60].Weight_n = Wgt_2_354;
         Mult_Buf[61].Feature_n = FeatureBuf_355;
         Mult_Buf[61].Weight_n = Wgt_2_355;
         Mult_Buf[62].Feature_n = FeatureBuf_356;
         Mult_Buf[62].Weight_n = Wgt_2_356;
         Mult_Buf[63].Feature_n = FeatureBuf_357;
         Mult_Buf[63].Weight_n = Wgt_2_357;
         Mult_Buf[64].Feature_n = FeatureBuf_358;
         Mult_Buf[64].Weight_n = Wgt_2_358;
         Mult_Buf[65].Feature_n = FeatureBuf_359;
         Mult_Buf[65].Weight_n = Wgt_2_359;
         Mult_Buf[66].Feature_n = FeatureBuf_360;
         Mult_Buf[66].Weight_n = Wgt_2_360;
         Mult_Buf[67].Feature_n = FeatureBuf_361;
         Mult_Buf[67].Weight_n = Wgt_2_361;
         Mult_Buf[68].Feature_n = FeatureBuf_362;
         Mult_Buf[68].Weight_n = Wgt_2_362;
         Mult_Buf[69].Feature_n = FeatureBuf_363;
         Mult_Buf[69].Weight_n = Wgt_2_363;
         Mult_Buf[70].Feature_n = FeatureBuf_364;
         Mult_Buf[70].Weight_n = Wgt_2_364;
         Mult_Buf[71].Feature_n = FeatureBuf_365;
         Mult_Buf[71].Weight_n = Wgt_2_365;
         Mult_Buf[72].Feature_n = FeatureBuf_366;
         Mult_Buf[72].Weight_n = Wgt_2_366;
         Mult_Buf[73].Feature_n = FeatureBuf_367;
         Mult_Buf[73].Weight_n = Wgt_2_367;
         Mult_Buf[74].Feature_n = FeatureBuf_368;
         Mult_Buf[74].Weight_n = Wgt_2_368;
         Mult_Buf[75].Feature_n = FeatureBuf_369;
         Mult_Buf[75].Weight_n = Wgt_2_369;
         Mult_Buf[76].Feature_n = FeatureBuf_370;
         Mult_Buf[76].Weight_n = Wgt_2_370;
         Mult_Buf[77].Feature_n = FeatureBuf_371;
         Mult_Buf[77].Weight_n = Wgt_2_371;
         Mult_Buf[78].Feature_n = FeatureBuf_372;
         Mult_Buf[78].Weight_n = Wgt_2_372;
         Mult_Buf[79].Feature_n = FeatureBuf_373;
         Mult_Buf[79].Weight_n = Wgt_2_373;
         Mult_Buf[80].Feature_n = FeatureBuf_374;
         Mult_Buf[80].Weight_n = Wgt_2_374;
         Mult_Buf[81].Feature_n = FeatureBuf_375;
         Mult_Buf[81].Weight_n = Wgt_2_375;
         Mult_Buf[82].Feature_n = FeatureBuf_376;
         Mult_Buf[82].Weight_n = Wgt_2_376;
         Mult_Buf[83].Feature_n = FeatureBuf_377;
         Mult_Buf[83].Weight_n = Wgt_2_377;
         Mult_Buf[84].Feature_n = FeatureBuf_378;
         Mult_Buf[84].Weight_n = Wgt_2_378;
         Mult_Buf[85].Feature_n = FeatureBuf_379;
         Mult_Buf[85].Weight_n = Wgt_2_379;
         Mult_Buf[86].Feature_n = FeatureBuf_380;
         Mult_Buf[86].Weight_n = Wgt_2_380;
         Mult_Buf[87].Feature_n = FeatureBuf_381;
         Mult_Buf[87].Weight_n = Wgt_2_381;
         Mult_Buf[88].Feature_n = FeatureBuf_382;
         Mult_Buf[88].Weight_n = Wgt_2_382;
         Mult_Buf[89].Feature_n = FeatureBuf_383;
         Mult_Buf[89].Weight_n = Wgt_2_383;
         Mult_Buf[90].Feature_n = FeatureBuf_384;
         Mult_Buf[90].Weight_n = Wgt_2_384;
         Mult_Buf[91].Feature_n = FeatureBuf_385;
         Mult_Buf[91].Weight_n = Wgt_2_385;
         Mult_Buf[92].Feature_n = FeatureBuf_386;
         Mult_Buf[92].Weight_n = Wgt_2_386;
         Mult_Buf[93].Feature_n = FeatureBuf_387;
         Mult_Buf[93].Weight_n = Wgt_2_387;
         Mult_Buf[94].Feature_n = FeatureBuf_388;
         Mult_Buf[94].Weight_n = Wgt_2_388;
         Mult_Buf[95].Feature_n = FeatureBuf_389;
         Mult_Buf[95].Weight_n = Wgt_2_389;
         Mult_Buf[96].Feature_n = FeatureBuf_390;
         Mult_Buf[96].Weight_n = Wgt_2_390;
         Mult_Buf[97].Feature_n = FeatureBuf_391;
         Mult_Buf[97].Weight_n = Wgt_2_391;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     end
    22:begin
     nxt_state = 23;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_392;
         Mult_Buf[0].Weight_n = Wgt_2_392;
         Mult_Buf[1].Feature_n = FeatureBuf_393;
         Mult_Buf[1].Weight_n = Wgt_2_393;
         Mult_Buf[2].Feature_n = FeatureBuf_394;
         Mult_Buf[2].Weight_n = Wgt_2_394;
         Mult_Buf[3].Feature_n = FeatureBuf_395;
         Mult_Buf[3].Weight_n = Wgt_2_395;
         Mult_Buf[4].Feature_n = FeatureBuf_396;
         Mult_Buf[4].Weight_n = Wgt_2_396;
         Mult_Buf[5].Feature_n = FeatureBuf_397;
         Mult_Buf[5].Weight_n = Wgt_2_397;
         Mult_Buf[6].Feature_n = FeatureBuf_398;
         Mult_Buf[6].Weight_n = Wgt_2_398;
         Mult_Buf[7].Feature_n = FeatureBuf_399;
         Mult_Buf[7].Weight_n = Wgt_2_399;
         Mult_Buf[8].Feature_n = FeatureBuf_400;
         Mult_Buf[8].Weight_n = Wgt_2_400;
         Mult_Buf[9].Feature_n = FeatureBuf_401;
         Mult_Buf[9].Weight_n = Wgt_2_401;
         Mult_Buf[10].Feature_n = FeatureBuf_402;
         Mult_Buf[10].Weight_n = Wgt_2_402;
         Mult_Buf[11].Feature_n = FeatureBuf_403;
         Mult_Buf[11].Weight_n = Wgt_2_403;
         Mult_Buf[12].Feature_n = FeatureBuf_404;
         Mult_Buf[12].Weight_n = Wgt_2_404;
         Mult_Buf[13].Feature_n = FeatureBuf_405;
         Mult_Buf[13].Weight_n = Wgt_2_405;
         Mult_Buf[14].Feature_n = FeatureBuf_406;
         Mult_Buf[14].Weight_n = Wgt_2_406;
         Mult_Buf[15].Feature_n = FeatureBuf_407;
         Mult_Buf[15].Weight_n = Wgt_2_407;
         Mult_Buf[16].Feature_n = FeatureBuf_408;
         Mult_Buf[16].Weight_n = Wgt_2_408;
         Mult_Buf[17].Feature_n = FeatureBuf_409;
         Mult_Buf[17].Weight_n = Wgt_2_409;
         Mult_Buf[18].Feature_n = FeatureBuf_410;
         Mult_Buf[18].Weight_n = Wgt_2_410;
         Mult_Buf[19].Feature_n = FeatureBuf_411;
         Mult_Buf[19].Weight_n = Wgt_2_411;
         Mult_Buf[20].Feature_n = FeatureBuf_412;
         Mult_Buf[20].Weight_n = Wgt_2_412;
         Mult_Buf[21].Feature_n = FeatureBuf_413;
         Mult_Buf[21].Weight_n = Wgt_2_413;
         Mult_Buf[22].Feature_n = FeatureBuf_414;
         Mult_Buf[22].Weight_n = Wgt_2_414;
         Mult_Buf[23].Feature_n = FeatureBuf_415;
         Mult_Buf[23].Weight_n = Wgt_2_415;
         Mult_Buf[24].Feature_n = FeatureBuf_416;
         Mult_Buf[24].Weight_n = Wgt_2_416;
         Mult_Buf[25].Feature_n = FeatureBuf_417;
         Mult_Buf[25].Weight_n = Wgt_2_417;
         Mult_Buf[26].Feature_n = FeatureBuf_418;
         Mult_Buf[26].Weight_n = Wgt_2_418;
         Mult_Buf[27].Feature_n = FeatureBuf_419;
         Mult_Buf[27].Weight_n = Wgt_2_419;
         Mult_Buf[28].Feature_n = FeatureBuf_420;
         Mult_Buf[28].Weight_n = Wgt_2_420;
         Mult_Buf[29].Feature_n = FeatureBuf_421;
         Mult_Buf[29].Weight_n = Wgt_2_421;
         Mult_Buf[30].Feature_n = FeatureBuf_422;
         Mult_Buf[30].Weight_n = Wgt_2_422;
         Mult_Buf[31].Feature_n = FeatureBuf_423;
         Mult_Buf[31].Weight_n = Wgt_2_423;
         Mult_Buf[32].Feature_n = FeatureBuf_424;
         Mult_Buf[32].Weight_n = Wgt_2_424;
         Mult_Buf[33].Feature_n = FeatureBuf_425;
         Mult_Buf[33].Weight_n = Wgt_2_425;
         Mult_Buf[34].Feature_n = FeatureBuf_426;
         Mult_Buf[34].Weight_n = Wgt_2_426;
         Mult_Buf[35].Feature_n = FeatureBuf_427;
         Mult_Buf[35].Weight_n = Wgt_2_427;
         Mult_Buf[36].Feature_n = FeatureBuf_428;
         Mult_Buf[36].Weight_n = Wgt_2_428;
         Mult_Buf[37].Feature_n = FeatureBuf_429;
         Mult_Buf[37].Weight_n = Wgt_2_429;
         Mult_Buf[38].Feature_n = FeatureBuf_430;
         Mult_Buf[38].Weight_n = Wgt_2_430;
         Mult_Buf[39].Feature_n = FeatureBuf_431;
         Mult_Buf[39].Weight_n = Wgt_2_431;
         Mult_Buf[40].Feature_n = FeatureBuf_432;
         Mult_Buf[40].Weight_n = Wgt_2_432;
         Mult_Buf[41].Feature_n = FeatureBuf_433;
         Mult_Buf[41].Weight_n = Wgt_2_433;
         Mult_Buf[42].Feature_n = FeatureBuf_434;
         Mult_Buf[42].Weight_n = Wgt_2_434;
         Mult_Buf[43].Feature_n = FeatureBuf_435;
         Mult_Buf[43].Weight_n = Wgt_2_435;
         Mult_Buf[44].Feature_n = FeatureBuf_436;
         Mult_Buf[44].Weight_n = Wgt_2_436;
         Mult_Buf[45].Feature_n = FeatureBuf_437;
         Mult_Buf[45].Weight_n = Wgt_2_437;
         Mult_Buf[46].Feature_n = FeatureBuf_438;
         Mult_Buf[46].Weight_n = Wgt_2_438;
         Mult_Buf[47].Feature_n = FeatureBuf_439;
         Mult_Buf[47].Weight_n = Wgt_2_439;
         Mult_Buf[48].Feature_n = FeatureBuf_440;
         Mult_Buf[48].Weight_n = Wgt_2_440;
         Mult_Buf[49].Feature_n = FeatureBuf_441;
         Mult_Buf[49].Weight_n = Wgt_2_441;
         Mult_Buf[50].Feature_n = FeatureBuf_442;
         Mult_Buf[50].Weight_n = Wgt_2_442;
         Mult_Buf[51].Feature_n = FeatureBuf_443;
         Mult_Buf[51].Weight_n = Wgt_2_443;
         Mult_Buf[52].Feature_n = FeatureBuf_444;
         Mult_Buf[52].Weight_n = Wgt_2_444;
         Mult_Buf[53].Feature_n = FeatureBuf_445;
         Mult_Buf[53].Weight_n = Wgt_2_445;
         Mult_Buf[54].Feature_n = FeatureBuf_446;
         Mult_Buf[54].Weight_n = Wgt_2_446;
         Mult_Buf[55].Feature_n = FeatureBuf_447;
         Mult_Buf[55].Weight_n = Wgt_2_447;
         Mult_Buf[56].Feature_n = FeatureBuf_448;
         Mult_Buf[56].Weight_n = Wgt_2_448;
         Mult_Buf[57].Feature_n = FeatureBuf_449;
         Mult_Buf[57].Weight_n = Wgt_2_449;
         Mult_Buf[58].Feature_n = FeatureBuf_450;
         Mult_Buf[58].Weight_n = Wgt_2_450;
         Mult_Buf[59].Feature_n = FeatureBuf_451;
         Mult_Buf[59].Weight_n = Wgt_2_451;
         Mult_Buf[60].Feature_n = FeatureBuf_452;
         Mult_Buf[60].Weight_n = Wgt_2_452;
         Mult_Buf[61].Feature_n = FeatureBuf_453;
         Mult_Buf[61].Weight_n = Wgt_2_453;
         Mult_Buf[62].Feature_n = FeatureBuf_454;
         Mult_Buf[62].Weight_n = Wgt_2_454;
         Mult_Buf[63].Feature_n = FeatureBuf_455;
         Mult_Buf[63].Weight_n = Wgt_2_455;
         Mult_Buf[64].Feature_n = FeatureBuf_456;
         Mult_Buf[64].Weight_n = Wgt_2_456;
         Mult_Buf[65].Feature_n = FeatureBuf_457;
         Mult_Buf[65].Weight_n = Wgt_2_457;
         Mult_Buf[66].Feature_n = FeatureBuf_458;
         Mult_Buf[66].Weight_n = Wgt_2_458;
         Mult_Buf[67].Feature_n = FeatureBuf_459;
         Mult_Buf[67].Weight_n = Wgt_2_459;
         Mult_Buf[68].Feature_n = FeatureBuf_460;
         Mult_Buf[68].Weight_n = Wgt_2_460;
         Mult_Buf[69].Feature_n = FeatureBuf_461;
         Mult_Buf[69].Weight_n = Wgt_2_461;
         Mult_Buf[70].Feature_n = FeatureBuf_462;
         Mult_Buf[70].Weight_n = Wgt_2_462;
         Mult_Buf[71].Feature_n = FeatureBuf_463;
         Mult_Buf[71].Weight_n = Wgt_2_463;
         Mult_Buf[72].Feature_n = FeatureBuf_464;
         Mult_Buf[72].Weight_n = Wgt_2_464;
         Mult_Buf[73].Feature_n = FeatureBuf_465;
         Mult_Buf[73].Weight_n = Wgt_2_465;
         Mult_Buf[74].Feature_n = FeatureBuf_466;
         Mult_Buf[74].Weight_n = Wgt_2_466;
         Mult_Buf[75].Feature_n = FeatureBuf_467;
         Mult_Buf[75].Weight_n = Wgt_2_467;
         Mult_Buf[76].Feature_n = FeatureBuf_468;
         Mult_Buf[76].Weight_n = Wgt_2_468;
         Mult_Buf[77].Feature_n = FeatureBuf_469;
         Mult_Buf[77].Weight_n = Wgt_2_469;
         Mult_Buf[78].Feature_n = FeatureBuf_470;
         Mult_Buf[78].Weight_n = Wgt_2_470;
         Mult_Buf[79].Feature_n = FeatureBuf_471;
         Mult_Buf[79].Weight_n = Wgt_2_471;
         Mult_Buf[80].Feature_n = FeatureBuf_472;
         Mult_Buf[80].Weight_n = Wgt_2_472;
         Mult_Buf[81].Feature_n = FeatureBuf_473;
         Mult_Buf[81].Weight_n = Wgt_2_473;
         Mult_Buf[82].Feature_n = FeatureBuf_474;
         Mult_Buf[82].Weight_n = Wgt_2_474;
         Mult_Buf[83].Feature_n = FeatureBuf_475;
         Mult_Buf[83].Weight_n = Wgt_2_475;
         Mult_Buf[84].Feature_n = FeatureBuf_476;
         Mult_Buf[84].Weight_n = Wgt_2_476;
         Mult_Buf[85].Feature_n = FeatureBuf_477;
         Mult_Buf[85].Weight_n = Wgt_2_477;
         Mult_Buf[86].Feature_n = FeatureBuf_478;
         Mult_Buf[86].Weight_n = Wgt_2_478;
         Mult_Buf[87].Feature_n = FeatureBuf_479;
         Mult_Buf[87].Weight_n = Wgt_2_479;
         Mult_Buf[88].Feature_n = FeatureBuf_480;
         Mult_Buf[88].Weight_n = Wgt_2_480;
         Mult_Buf[89].Feature_n = FeatureBuf_481;
         Mult_Buf[89].Weight_n = Wgt_2_481;
         Mult_Buf[90].Feature_n = FeatureBuf_482;
         Mult_Buf[90].Weight_n = Wgt_2_482;
         Mult_Buf[91].Feature_n = FeatureBuf_483;
         Mult_Buf[91].Weight_n = Wgt_2_483;
         Mult_Buf[92].Feature_n = FeatureBuf_484;
         Mult_Buf[92].Weight_n = Wgt_2_484;
         Mult_Buf[93].Feature_n = FeatureBuf_485;
         Mult_Buf[93].Weight_n = Wgt_2_485;
         Mult_Buf[94].Feature_n = FeatureBuf_486;
         Mult_Buf[94].Weight_n = Wgt_2_486;
         Mult_Buf[95].Feature_n = FeatureBuf_487;
         Mult_Buf[95].Weight_n = Wgt_2_487;
         Mult_Buf[96].Feature_n = FeatureBuf_488;
         Mult_Buf[96].Weight_n = Wgt_2_488;
         Mult_Buf[97].Feature_n = FeatureBuf_489;
         Mult_Buf[97].Weight_n = Wgt_2_489;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     end
    23:begin
     nxt_state = 24;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_490;
         Mult_Buf[0].Weight_n = Wgt_2_490;
         Mult_Buf[1].Feature_n = FeatureBuf_491;
         Mult_Buf[1].Weight_n = Wgt_2_491;
         Mult_Buf[2].Feature_n = FeatureBuf_492;
         Mult_Buf[2].Weight_n = Wgt_2_492;
         Mult_Buf[3].Feature_n = FeatureBuf_493;
         Mult_Buf[3].Weight_n = Wgt_2_493;
         Mult_Buf[4].Feature_n = FeatureBuf_494;
         Mult_Buf[4].Weight_n = Wgt_2_494;
         Mult_Buf[5].Feature_n = FeatureBuf_495;
         Mult_Buf[5].Weight_n = Wgt_2_495;
         Mult_Buf[6].Feature_n = FeatureBuf_496;
         Mult_Buf[6].Weight_n = Wgt_2_496;
         Mult_Buf[7].Feature_n = FeatureBuf_497;
         Mult_Buf[7].Weight_n = Wgt_2_497;
         Mult_Buf[8].Feature_n = FeatureBuf_498;
         Mult_Buf[8].Weight_n = Wgt_2_498;
         Mult_Buf[9].Feature_n = FeatureBuf_499;
         Mult_Buf[9].Weight_n = Wgt_2_499;
         Mult_Buf[10].Feature_n = FeatureBuf_500;
         Mult_Buf[10].Weight_n = Wgt_2_500;
         Mult_Buf[11].Feature_n = FeatureBuf_501;
         Mult_Buf[11].Weight_n = Wgt_2_501;
         Mult_Buf[12].Feature_n = FeatureBuf_502;
         Mult_Buf[12].Weight_n = Wgt_2_502;
         Mult_Buf[13].Feature_n = FeatureBuf_503;
         Mult_Buf[13].Weight_n = Wgt_2_503;
         Mult_Buf[14].Feature_n = FeatureBuf_504;
         Mult_Buf[14].Weight_n = Wgt_2_504;
         Mult_Buf[15].Feature_n = FeatureBuf_505;
         Mult_Buf[15].Weight_n = Wgt_2_505;
         Mult_Buf[16].Feature_n = FeatureBuf_506;
         Mult_Buf[16].Weight_n = Wgt_2_506;
         Mult_Buf[17].Feature_n = FeatureBuf_507;
         Mult_Buf[17].Weight_n = Wgt_2_507;
         Mult_Buf[18].Feature_n = FeatureBuf_508;
         Mult_Buf[18].Weight_n = Wgt_2_508;
         Mult_Buf[19].Feature_n = FeatureBuf_509;
         Mult_Buf[19].Weight_n = Wgt_2_509;
         Mult_Buf[20].Feature_n = FeatureBuf_510;
         Mult_Buf[20].Weight_n = Wgt_2_510;
         Mult_Buf[21].Feature_n = FeatureBuf_511;
         Mult_Buf[21].Weight_n = Wgt_2_511;
         Mult_Buf[22].Feature_n = FeatureBuf_512;
         Mult_Buf[22].Weight_n = Wgt_2_512;
         Mult_Buf[23].Feature_n = FeatureBuf_513;
         Mult_Buf[23].Weight_n = Wgt_2_513;
         Mult_Buf[24].Feature_n = FeatureBuf_514;
         Mult_Buf[24].Weight_n = Wgt_2_514;
         Mult_Buf[25].Feature_n = FeatureBuf_515;
         Mult_Buf[25].Weight_n = Wgt_2_515;
         Mult_Buf[26].Feature_n = FeatureBuf_516;
         Mult_Buf[26].Weight_n = Wgt_2_516;
         Mult_Buf[27].Feature_n = FeatureBuf_517;
         Mult_Buf[27].Weight_n = Wgt_2_517;
         Mult_Buf[28].Feature_n = FeatureBuf_518;
         Mult_Buf[28].Weight_n = Wgt_2_518;
         Mult_Buf[29].Feature_n = FeatureBuf_519;
         Mult_Buf[29].Weight_n = Wgt_2_519;
         Mult_Buf[30].Feature_n = FeatureBuf_520;
         Mult_Buf[30].Weight_n = Wgt_2_520;
         Mult_Buf[31].Feature_n = FeatureBuf_521;
         Mult_Buf[31].Weight_n = Wgt_2_521;
         Mult_Buf[32].Feature_n = FeatureBuf_522;
         Mult_Buf[32].Weight_n = Wgt_2_522;
         Mult_Buf[33].Feature_n = FeatureBuf_523;
         Mult_Buf[33].Weight_n = Wgt_2_523;
         Mult_Buf[34].Feature_n = FeatureBuf_524;
         Mult_Buf[34].Weight_n = Wgt_2_524;
         Mult_Buf[35].Feature_n = FeatureBuf_525;
         Mult_Buf[35].Weight_n = Wgt_2_525;
         Mult_Buf[36].Feature_n = FeatureBuf_526;
         Mult_Buf[36].Weight_n = Wgt_2_526;
         Mult_Buf[37].Feature_n = FeatureBuf_527;
         Mult_Buf[37].Weight_n = Wgt_2_527;
         Mult_Buf[38].Feature_n = FeatureBuf_528;
         Mult_Buf[38].Weight_n = Wgt_2_528;
         Mult_Buf[39].Feature_n = FeatureBuf_529;
         Mult_Buf[39].Weight_n = Wgt_2_529;
         Mult_Buf[40].Feature_n = FeatureBuf_530;
         Mult_Buf[40].Weight_n = Wgt_2_530;
         Mult_Buf[41].Feature_n = FeatureBuf_531;
         Mult_Buf[41].Weight_n = Wgt_2_531;
         Mult_Buf[42].Feature_n = FeatureBuf_532;
         Mult_Buf[42].Weight_n = Wgt_2_532;
         Mult_Buf[43].Feature_n = FeatureBuf_533;
         Mult_Buf[43].Weight_n = Wgt_2_533;
         Mult_Buf[44].Feature_n = FeatureBuf_534;
         Mult_Buf[44].Weight_n = Wgt_2_534;
         Mult_Buf[45].Feature_n = FeatureBuf_535;
         Mult_Buf[45].Weight_n = Wgt_2_535;
         Mult_Buf[46].Feature_n = FeatureBuf_536;
         Mult_Buf[46].Weight_n = Wgt_2_536;
         Mult_Buf[47].Feature_n = FeatureBuf_537;
         Mult_Buf[47].Weight_n = Wgt_2_537;
         Mult_Buf[48].Feature_n = FeatureBuf_538;
         Mult_Buf[48].Weight_n = Wgt_2_538;
         Mult_Buf[49].Feature_n = FeatureBuf_539;
         Mult_Buf[49].Weight_n = Wgt_2_539;
         Mult_Buf[50].Feature_n = FeatureBuf_540;
         Mult_Buf[50].Weight_n = Wgt_2_540;
         Mult_Buf[51].Feature_n = FeatureBuf_541;
         Mult_Buf[51].Weight_n = Wgt_2_541;
         Mult_Buf[52].Feature_n = FeatureBuf_542;
         Mult_Buf[52].Weight_n = Wgt_2_542;
         Mult_Buf[53].Feature_n = FeatureBuf_543;
         Mult_Buf[53].Weight_n = Wgt_2_543;
         Mult_Buf[54].Feature_n = FeatureBuf_544;
         Mult_Buf[54].Weight_n = Wgt_2_544;
         Mult_Buf[55].Feature_n = FeatureBuf_545;
         Mult_Buf[55].Weight_n = Wgt_2_545;
         Mult_Buf[56].Feature_n = FeatureBuf_546;
         Mult_Buf[56].Weight_n = Wgt_2_546;
         Mult_Buf[57].Feature_n = FeatureBuf_547;
         Mult_Buf[57].Weight_n = Wgt_2_547;
         Mult_Buf[58].Feature_n = FeatureBuf_548;
         Mult_Buf[58].Weight_n = Wgt_2_548;
         Mult_Buf[59].Feature_n = FeatureBuf_549;
         Mult_Buf[59].Weight_n = Wgt_2_549;
         Mult_Buf[60].Feature_n = FeatureBuf_550;
         Mult_Buf[60].Weight_n = Wgt_2_550;
         Mult_Buf[61].Feature_n = FeatureBuf_551;
         Mult_Buf[61].Weight_n = Wgt_2_551;
         Mult_Buf[62].Feature_n = FeatureBuf_552;
         Mult_Buf[62].Weight_n = Wgt_2_552;
         Mult_Buf[63].Feature_n = FeatureBuf_553;
         Mult_Buf[63].Weight_n = Wgt_2_553;
         Mult_Buf[64].Feature_n = FeatureBuf_554;
         Mult_Buf[64].Weight_n = Wgt_2_554;
         Mult_Buf[65].Feature_n = FeatureBuf_555;
         Mult_Buf[65].Weight_n = Wgt_2_555;
         Mult_Buf[66].Feature_n = FeatureBuf_556;
         Mult_Buf[66].Weight_n = Wgt_2_556;
         Mult_Buf[67].Feature_n = FeatureBuf_557;
         Mult_Buf[67].Weight_n = Wgt_2_557;
         Mult_Buf[68].Feature_n = FeatureBuf_558;
         Mult_Buf[68].Weight_n = Wgt_2_558;
         Mult_Buf[69].Feature_n = FeatureBuf_559;
         Mult_Buf[69].Weight_n = Wgt_2_559;
         Mult_Buf[70].Feature_n = FeatureBuf_560;
         Mult_Buf[70].Weight_n = Wgt_2_560;
         Mult_Buf[71].Feature_n = FeatureBuf_561;
         Mult_Buf[71].Weight_n = Wgt_2_561;
         Mult_Buf[72].Feature_n = FeatureBuf_562;
         Mult_Buf[72].Weight_n = Wgt_2_562;
         Mult_Buf[73].Feature_n = FeatureBuf_563;
         Mult_Buf[73].Weight_n = Wgt_2_563;
         Mult_Buf[74].Feature_n = FeatureBuf_564;
         Mult_Buf[74].Weight_n = Wgt_2_564;
         Mult_Buf[75].Feature_n = FeatureBuf_565;
         Mult_Buf[75].Weight_n = Wgt_2_565;
         Mult_Buf[76].Feature_n = FeatureBuf_566;
         Mult_Buf[76].Weight_n = Wgt_2_566;
         Mult_Buf[77].Feature_n = FeatureBuf_567;
         Mult_Buf[77].Weight_n = Wgt_2_567;
         Mult_Buf[78].Feature_n = FeatureBuf_568;
         Mult_Buf[78].Weight_n = Wgt_2_568;
         Mult_Buf[79].Feature_n = FeatureBuf_569;
         Mult_Buf[79].Weight_n = Wgt_2_569;
         Mult_Buf[80].Feature_n = FeatureBuf_570;
         Mult_Buf[80].Weight_n = Wgt_2_570;
         Mult_Buf[81].Feature_n = FeatureBuf_571;
         Mult_Buf[81].Weight_n = Wgt_2_571;
         Mult_Buf[82].Feature_n = FeatureBuf_572;
         Mult_Buf[82].Weight_n = Wgt_2_572;
         Mult_Buf[83].Feature_n = FeatureBuf_573;
         Mult_Buf[83].Weight_n = Wgt_2_573;
         Mult_Buf[84].Feature_n = FeatureBuf_574;
         Mult_Buf[84].Weight_n = Wgt_2_574;
         Mult_Buf[85].Feature_n = FeatureBuf_575;
         Mult_Buf[85].Weight_n = Wgt_2_575;
         Mult_Buf[86].Feature_n = FeatureBuf_576;
         Mult_Buf[86].Weight_n = Wgt_2_576;
         Mult_Buf[87].Feature_n = FeatureBuf_577;
         Mult_Buf[87].Weight_n = Wgt_2_577;
         Mult_Buf[88].Feature_n = FeatureBuf_578;
         Mult_Buf[88].Weight_n = Wgt_2_578;
         Mult_Buf[89].Feature_n = FeatureBuf_579;
         Mult_Buf[89].Weight_n = Wgt_2_579;
         Mult_Buf[90].Feature_n = FeatureBuf_580;
         Mult_Buf[90].Weight_n = Wgt_2_580;
         Mult_Buf[91].Feature_n = FeatureBuf_581;
         Mult_Buf[91].Weight_n = Wgt_2_581;
         Mult_Buf[92].Feature_n = FeatureBuf_582;
         Mult_Buf[92].Weight_n = Wgt_2_582;
         Mult_Buf[93].Feature_n = FeatureBuf_583;
         Mult_Buf[93].Weight_n = Wgt_2_583;
         Mult_Buf[94].Feature_n = FeatureBuf_584;
         Mult_Buf[94].Weight_n = Wgt_2_584;
         Mult_Buf[95].Feature_n = FeatureBuf_585;
         Mult_Buf[95].Weight_n = Wgt_2_585;
         Mult_Buf[96].Feature_n = FeatureBuf_586;
         Mult_Buf[96].Weight_n = Wgt_2_586;
         Mult_Buf[97].Feature_n = FeatureBuf_587;
         Mult_Buf[97].Weight_n = Wgt_2_587;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     end
    24:begin
     nxt_state = 25;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_588;
         Mult_Buf[0].Weight_n = Wgt_2_588;
         Mult_Buf[1].Feature_n = FeatureBuf_589;
         Mult_Buf[1].Weight_n = Wgt_2_589;
         Mult_Buf[2].Feature_n = FeatureBuf_590;
         Mult_Buf[2].Weight_n = Wgt_2_590;
         Mult_Buf[3].Feature_n = FeatureBuf_591;
         Mult_Buf[3].Weight_n = Wgt_2_591;
         Mult_Buf[4].Feature_n = FeatureBuf_592;
         Mult_Buf[4].Weight_n = Wgt_2_592;
         Mult_Buf[5].Feature_n = FeatureBuf_593;
         Mult_Buf[5].Weight_n = Wgt_2_593;
         Mult_Buf[6].Feature_n = FeatureBuf_594;
         Mult_Buf[6].Weight_n = Wgt_2_594;
         Mult_Buf[7].Feature_n = FeatureBuf_595;
         Mult_Buf[7].Weight_n = Wgt_2_595;
         Mult_Buf[8].Feature_n = FeatureBuf_596;
         Mult_Buf[8].Weight_n = Wgt_2_596;
         Mult_Buf[9].Feature_n = FeatureBuf_597;
         Mult_Buf[9].Weight_n = Wgt_2_597;
         Mult_Buf[10].Feature_n = FeatureBuf_598;
         Mult_Buf[10].Weight_n = Wgt_2_598;
         Mult_Buf[11].Feature_n = FeatureBuf_599;
         Mult_Buf[11].Weight_n = Wgt_2_599;
         Mult_Buf[12].Feature_n = FeatureBuf_600;
         Mult_Buf[12].Weight_n = Wgt_2_600;
         Mult_Buf[13].Feature_n = FeatureBuf_601;
         Mult_Buf[13].Weight_n = Wgt_2_601;
         Mult_Buf[14].Feature_n = FeatureBuf_602;
         Mult_Buf[14].Weight_n = Wgt_2_602;
         Mult_Buf[15].Feature_n = FeatureBuf_603;
         Mult_Buf[15].Weight_n = Wgt_2_603;
         Mult_Buf[16].Feature_n = FeatureBuf_604;
         Mult_Buf[16].Weight_n = Wgt_2_604;
         Mult_Buf[17].Feature_n = FeatureBuf_605;
         Mult_Buf[17].Weight_n = Wgt_2_605;
         Mult_Buf[18].Feature_n = FeatureBuf_606;
         Mult_Buf[18].Weight_n = Wgt_2_606;
         Mult_Buf[19].Feature_n = FeatureBuf_607;
         Mult_Buf[19].Weight_n = Wgt_2_607;
         Mult_Buf[20].Feature_n = FeatureBuf_608;
         Mult_Buf[20].Weight_n = Wgt_2_608;
         Mult_Buf[21].Feature_n = FeatureBuf_609;
         Mult_Buf[21].Weight_n = Wgt_2_609;
         Mult_Buf[22].Feature_n = FeatureBuf_610;
         Mult_Buf[22].Weight_n = Wgt_2_610;
         Mult_Buf[23].Feature_n = FeatureBuf_611;
         Mult_Buf[23].Weight_n = Wgt_2_611;
         Mult_Buf[24].Feature_n = FeatureBuf_612;
         Mult_Buf[24].Weight_n = Wgt_2_612;
         Mult_Buf[25].Feature_n = FeatureBuf_613;
         Mult_Buf[25].Weight_n = Wgt_2_613;
         Mult_Buf[26].Feature_n = FeatureBuf_614;
         Mult_Buf[26].Weight_n = Wgt_2_614;
         Mult_Buf[27].Feature_n = FeatureBuf_615;
         Mult_Buf[27].Weight_n = Wgt_2_615;
         Mult_Buf[28].Feature_n = FeatureBuf_616;
         Mult_Buf[28].Weight_n = Wgt_2_616;
         Mult_Buf[29].Feature_n = FeatureBuf_617;
         Mult_Buf[29].Weight_n = Wgt_2_617;
         Mult_Buf[30].Feature_n = FeatureBuf_618;
         Mult_Buf[30].Weight_n = Wgt_2_618;
         Mult_Buf[31].Feature_n = FeatureBuf_619;
         Mult_Buf[31].Weight_n = Wgt_2_619;
         Mult_Buf[32].Feature_n = FeatureBuf_620;
         Mult_Buf[32].Weight_n = Wgt_2_620;
         Mult_Buf[33].Feature_n = FeatureBuf_621;
         Mult_Buf[33].Weight_n = Wgt_2_621;
         Mult_Buf[34].Feature_n = FeatureBuf_622;
         Mult_Buf[34].Weight_n = Wgt_2_622;
         Mult_Buf[35].Feature_n = FeatureBuf_623;
         Mult_Buf[35].Weight_n = Wgt_2_623;
         Mult_Buf[36].Feature_n = FeatureBuf_624;
         Mult_Buf[36].Weight_n = Wgt_2_624;
         Mult_Buf[37].Feature_n = FeatureBuf_625;
         Mult_Buf[37].Weight_n = Wgt_2_625;
         Mult_Buf[38].Feature_n = FeatureBuf_626;
         Mult_Buf[38].Weight_n = Wgt_2_626;
         Mult_Buf[39].Feature_n = FeatureBuf_627;
         Mult_Buf[39].Weight_n = Wgt_2_627;
         Mult_Buf[40].Feature_n = FeatureBuf_628;
         Mult_Buf[40].Weight_n = Wgt_2_628;
         Mult_Buf[41].Feature_n = FeatureBuf_629;
         Mult_Buf[41].Weight_n = Wgt_2_629;
         Mult_Buf[42].Feature_n = FeatureBuf_630;
         Mult_Buf[42].Weight_n = Wgt_2_630;
         Mult_Buf[43].Feature_n = FeatureBuf_631;
         Mult_Buf[43].Weight_n = Wgt_2_631;
         Mult_Buf[44].Feature_n = FeatureBuf_632;
         Mult_Buf[44].Weight_n = Wgt_2_632;
         Mult_Buf[45].Feature_n = FeatureBuf_633;
         Mult_Buf[45].Weight_n = Wgt_2_633;
         Mult_Buf[46].Feature_n = FeatureBuf_634;
         Mult_Buf[46].Weight_n = Wgt_2_634;
         Mult_Buf[47].Feature_n = FeatureBuf_635;
         Mult_Buf[47].Weight_n = Wgt_2_635;
         Mult_Buf[48].Feature_n = FeatureBuf_636;
         Mult_Buf[48].Weight_n = Wgt_2_636;
         Mult_Buf[49].Feature_n = FeatureBuf_637;
         Mult_Buf[49].Weight_n = Wgt_2_637;
         Mult_Buf[50].Feature_n = FeatureBuf_638;
         Mult_Buf[50].Weight_n = Wgt_2_638;
         Mult_Buf[51].Feature_n = FeatureBuf_639;
         Mult_Buf[51].Weight_n = Wgt_2_639;
         Mult_Buf[52].Feature_n = FeatureBuf_640;
         Mult_Buf[52].Weight_n = Wgt_2_640;
         Mult_Buf[53].Feature_n = FeatureBuf_641;
         Mult_Buf[53].Weight_n = Wgt_2_641;
         Mult_Buf[54].Feature_n = FeatureBuf_642;
         Mult_Buf[54].Weight_n = Wgt_2_642;
         Mult_Buf[55].Feature_n = FeatureBuf_643;
         Mult_Buf[55].Weight_n = Wgt_2_643;
         Mult_Buf[56].Feature_n = FeatureBuf_644;
         Mult_Buf[56].Weight_n = Wgt_2_644;
         Mult_Buf[57].Feature_n = FeatureBuf_645;
         Mult_Buf[57].Weight_n = Wgt_2_645;
         Mult_Buf[58].Feature_n = FeatureBuf_646;
         Mult_Buf[58].Weight_n = Wgt_2_646;
         Mult_Buf[59].Feature_n = FeatureBuf_647;
         Mult_Buf[59].Weight_n = Wgt_2_647;
         Mult_Buf[60].Feature_n = FeatureBuf_648;
         Mult_Buf[60].Weight_n = Wgt_2_648;
         Mult_Buf[61].Feature_n = FeatureBuf_649;
         Mult_Buf[61].Weight_n = Wgt_2_649;
         Mult_Buf[62].Feature_n = FeatureBuf_650;
         Mult_Buf[62].Weight_n = Wgt_2_650;
         Mult_Buf[63].Feature_n = FeatureBuf_651;
         Mult_Buf[63].Weight_n = Wgt_2_651;
         Mult_Buf[64].Feature_n = FeatureBuf_652;
         Mult_Buf[64].Weight_n = Wgt_2_652;
         Mult_Buf[65].Feature_n = FeatureBuf_653;
         Mult_Buf[65].Weight_n = Wgt_2_653;
         Mult_Buf[66].Feature_n = FeatureBuf_654;
         Mult_Buf[66].Weight_n = Wgt_2_654;
         Mult_Buf[67].Feature_n = FeatureBuf_655;
         Mult_Buf[67].Weight_n = Wgt_2_655;
         Mult_Buf[68].Feature_n = FeatureBuf_656;
         Mult_Buf[68].Weight_n = Wgt_2_656;
         Mult_Buf[69].Feature_n = FeatureBuf_657;
         Mult_Buf[69].Weight_n = Wgt_2_657;
         Mult_Buf[70].Feature_n = FeatureBuf_658;
         Mult_Buf[70].Weight_n = Wgt_2_658;
         Mult_Buf[71].Feature_n = FeatureBuf_659;
         Mult_Buf[71].Weight_n = Wgt_2_659;
         Mult_Buf[72].Feature_n = FeatureBuf_660;
         Mult_Buf[72].Weight_n = Wgt_2_660;
         Mult_Buf[73].Feature_n = FeatureBuf_661;
         Mult_Buf[73].Weight_n = Wgt_2_661;
         Mult_Buf[74].Feature_n = FeatureBuf_662;
         Mult_Buf[74].Weight_n = Wgt_2_662;
         Mult_Buf[75].Feature_n = FeatureBuf_663;
         Mult_Buf[75].Weight_n = Wgt_2_663;
         Mult_Buf[76].Feature_n = FeatureBuf_664;
         Mult_Buf[76].Weight_n = Wgt_2_664;
         Mult_Buf[77].Feature_n = FeatureBuf_665;
         Mult_Buf[77].Weight_n = Wgt_2_665;
         Mult_Buf[78].Feature_n = FeatureBuf_666;
         Mult_Buf[78].Weight_n = Wgt_2_666;
         Mult_Buf[79].Feature_n = FeatureBuf_667;
         Mult_Buf[79].Weight_n = Wgt_2_667;
         Mult_Buf[80].Feature_n = FeatureBuf_668;
         Mult_Buf[80].Weight_n = Wgt_2_668;
         Mult_Buf[81].Feature_n = FeatureBuf_669;
         Mult_Buf[81].Weight_n = Wgt_2_669;
         Mult_Buf[82].Feature_n = FeatureBuf_670;
         Mult_Buf[82].Weight_n = Wgt_2_670;
         Mult_Buf[83].Feature_n = FeatureBuf_671;
         Mult_Buf[83].Weight_n = Wgt_2_671;
         Mult_Buf[84].Feature_n = FeatureBuf_672;
         Mult_Buf[84].Weight_n = Wgt_2_672;
         Mult_Buf[85].Feature_n = FeatureBuf_673;
         Mult_Buf[85].Weight_n = Wgt_2_673;
         Mult_Buf[86].Feature_n = FeatureBuf_674;
         Mult_Buf[86].Weight_n = Wgt_2_674;
         Mult_Buf[87].Feature_n = FeatureBuf_675;
         Mult_Buf[87].Weight_n = Wgt_2_675;
         Mult_Buf[88].Feature_n = FeatureBuf_676;
         Mult_Buf[88].Weight_n = Wgt_2_676;
         Mult_Buf[89].Feature_n = FeatureBuf_677;
         Mult_Buf[89].Weight_n = Wgt_2_677;
         Mult_Buf[90].Feature_n = FeatureBuf_678;
         Mult_Buf[90].Weight_n = Wgt_2_678;
         Mult_Buf[91].Feature_n = FeatureBuf_679;
         Mult_Buf[91].Weight_n = Wgt_2_679;
         Mult_Buf[92].Feature_n = FeatureBuf_680;
         Mult_Buf[92].Weight_n = Wgt_2_680;
         Mult_Buf[93].Feature_n = FeatureBuf_681;
         Mult_Buf[93].Weight_n = Wgt_2_681;
         Mult_Buf[94].Feature_n = FeatureBuf_682;
         Mult_Buf[94].Weight_n = Wgt_2_682;
         Mult_Buf[95].Feature_n = FeatureBuf_683;
         Mult_Buf[95].Weight_n = Wgt_2_683;
         Mult_Buf[96].Feature_n = FeatureBuf_684;
         Mult_Buf[96].Weight_n = Wgt_2_684;
         Mult_Buf[97].Feature_n = FeatureBuf_685;
         Mult_Buf[97].Weight_n = Wgt_2_685;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     //Collect Partial result form Adder
         Res_0_0_n = Part_Res;
     end
    25:begin
     nxt_state = 26;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_686;
         Mult_Buf[0].Weight_n = Wgt_2_686;
         Mult_Buf[1].Feature_n = FeatureBuf_687;
         Mult_Buf[1].Weight_n = Wgt_2_687;
         Mult_Buf[2].Feature_n = FeatureBuf_688;
         Mult_Buf[2].Weight_n = Wgt_2_688;
         Mult_Buf[3].Feature_n = FeatureBuf_689;
         Mult_Buf[3].Weight_n = Wgt_2_689;
         Mult_Buf[4].Feature_n = FeatureBuf_690;
         Mult_Buf[4].Weight_n = Wgt_2_690;
         Mult_Buf[5].Feature_n = FeatureBuf_691;
         Mult_Buf[5].Weight_n = Wgt_2_691;
         Mult_Buf[6].Feature_n = FeatureBuf_692;
         Mult_Buf[6].Weight_n = Wgt_2_692;
         Mult_Buf[7].Feature_n = FeatureBuf_693;
         Mult_Buf[7].Weight_n = Wgt_2_693;
         Mult_Buf[8].Feature_n = FeatureBuf_694;
         Mult_Buf[8].Weight_n = Wgt_2_694;
         Mult_Buf[9].Feature_n = FeatureBuf_695;
         Mult_Buf[9].Weight_n = Wgt_2_695;
         Mult_Buf[10].Feature_n = FeatureBuf_696;
         Mult_Buf[10].Weight_n = Wgt_2_696;
         Mult_Buf[11].Feature_n = FeatureBuf_697;
         Mult_Buf[11].Weight_n = Wgt_2_697;
         Mult_Buf[12].Feature_n = FeatureBuf_698;
         Mult_Buf[12].Weight_n = Wgt_2_698;
         Mult_Buf[13].Feature_n = FeatureBuf_699;
         Mult_Buf[13].Weight_n = Wgt_2_699;
         Mult_Buf[14].Feature_n = FeatureBuf_700;
         Mult_Buf[14].Weight_n = Wgt_2_700;
         Mult_Buf[15].Feature_n = FeatureBuf_701;
         Mult_Buf[15].Weight_n = Wgt_2_701;
         Mult_Buf[16].Feature_n = FeatureBuf_702;
         Mult_Buf[16].Weight_n = Wgt_2_702;
         Mult_Buf[17].Feature_n = FeatureBuf_703;
         Mult_Buf[17].Weight_n = Wgt_2_703;
         Mult_Buf[18].Feature_n = FeatureBuf_704;
         Mult_Buf[18].Weight_n = Wgt_2_704;
         Mult_Buf[19].Feature_n = FeatureBuf_705;
         Mult_Buf[19].Weight_n = Wgt_2_705;
         Mult_Buf[20].Feature_n = FeatureBuf_706;
         Mult_Buf[20].Weight_n = Wgt_2_706;
         Mult_Buf[21].Feature_n = FeatureBuf_707;
         Mult_Buf[21].Weight_n = Wgt_2_707;
         Mult_Buf[22].Feature_n = FeatureBuf_708;
         Mult_Buf[22].Weight_n = Wgt_2_708;
         Mult_Buf[23].Feature_n = FeatureBuf_709;
         Mult_Buf[23].Weight_n = Wgt_2_709;
         Mult_Buf[24].Feature_n = FeatureBuf_710;
         Mult_Buf[24].Weight_n = Wgt_2_710;
         Mult_Buf[25].Feature_n = FeatureBuf_711;
         Mult_Buf[25].Weight_n = Wgt_2_711;
         Mult_Buf[26].Feature_n = FeatureBuf_712;
         Mult_Buf[26].Weight_n = Wgt_2_712;
         Mult_Buf[27].Feature_n = FeatureBuf_713;
         Mult_Buf[27].Weight_n = Wgt_2_713;
         Mult_Buf[28].Feature_n = FeatureBuf_714;
         Mult_Buf[28].Weight_n = Wgt_2_714;
         Mult_Buf[29].Feature_n = FeatureBuf_715;
         Mult_Buf[29].Weight_n = Wgt_2_715;
         Mult_Buf[30].Feature_n = FeatureBuf_716;
         Mult_Buf[30].Weight_n = Wgt_2_716;
         Mult_Buf[31].Feature_n = FeatureBuf_717;
         Mult_Buf[31].Weight_n = Wgt_2_717;
         Mult_Buf[32].Feature_n = FeatureBuf_718;
         Mult_Buf[32].Weight_n = Wgt_2_718;
         Mult_Buf[33].Feature_n = FeatureBuf_719;
         Mult_Buf[33].Weight_n = Wgt_2_719;
         Mult_Buf[34].Feature_n = FeatureBuf_720;
         Mult_Buf[34].Weight_n = Wgt_2_720;
         Mult_Buf[35].Feature_n = FeatureBuf_721;
         Mult_Buf[35].Weight_n = Wgt_2_721;
         Mult_Buf[36].Feature_n = FeatureBuf_722;
         Mult_Buf[36].Weight_n = Wgt_2_722;
         Mult_Buf[37].Feature_n = FeatureBuf_723;
         Mult_Buf[37].Weight_n = Wgt_2_723;
         Mult_Buf[38].Feature_n = FeatureBuf_724;
         Mult_Buf[38].Weight_n = Wgt_2_724;
         Mult_Buf[39].Feature_n = FeatureBuf_725;
         Mult_Buf[39].Weight_n = Wgt_2_725;
         Mult_Buf[40].Feature_n = FeatureBuf_726;
         Mult_Buf[40].Weight_n = Wgt_2_726;
         Mult_Buf[41].Feature_n = FeatureBuf_727;
         Mult_Buf[41].Weight_n = Wgt_2_727;
         Mult_Buf[42].Feature_n = FeatureBuf_728;
         Mult_Buf[42].Weight_n = Wgt_2_728;
         Mult_Buf[43].Feature_n = FeatureBuf_729;
         Mult_Buf[43].Weight_n = Wgt_2_729;
         Mult_Buf[44].Feature_n = FeatureBuf_730;
         Mult_Buf[44].Weight_n = Wgt_2_730;
         Mult_Buf[45].Feature_n = FeatureBuf_731;
         Mult_Buf[45].Weight_n = Wgt_2_731;
         Mult_Buf[46].Feature_n = FeatureBuf_732;
         Mult_Buf[46].Weight_n = Wgt_2_732;
         Mult_Buf[47].Feature_n = FeatureBuf_733;
         Mult_Buf[47].Weight_n = Wgt_2_733;
         Mult_Buf[48].Feature_n = FeatureBuf_734;
         Mult_Buf[48].Weight_n = Wgt_2_734;
         Mult_Buf[49].Feature_n = FeatureBuf_735;
         Mult_Buf[49].Weight_n = Wgt_2_735;
         Mult_Buf[50].Feature_n = FeatureBuf_736;
         Mult_Buf[50].Weight_n = Wgt_2_736;
         Mult_Buf[51].Feature_n = FeatureBuf_737;
         Mult_Buf[51].Weight_n = Wgt_2_737;
         Mult_Buf[52].Feature_n = FeatureBuf_738;
         Mult_Buf[52].Weight_n = Wgt_2_738;
         Mult_Buf[53].Feature_n = FeatureBuf_739;
         Mult_Buf[53].Weight_n = Wgt_2_739;
         Mult_Buf[54].Feature_n = FeatureBuf_740;
         Mult_Buf[54].Weight_n = Wgt_2_740;
         Mult_Buf[55].Feature_n = FeatureBuf_741;
         Mult_Buf[55].Weight_n = Wgt_2_741;
         Mult_Buf[56].Feature_n = FeatureBuf_742;
         Mult_Buf[56].Weight_n = Wgt_2_742;
         Mult_Buf[57].Feature_n = FeatureBuf_743;
         Mult_Buf[57].Weight_n = Wgt_2_743;
         Mult_Buf[58].Feature_n = FeatureBuf_744;
         Mult_Buf[58].Weight_n = Wgt_2_744;
         Mult_Buf[59].Feature_n = FeatureBuf_745;
         Mult_Buf[59].Weight_n = Wgt_2_745;
         Mult_Buf[60].Feature_n = FeatureBuf_746;
         Mult_Buf[60].Weight_n = Wgt_2_746;
         Mult_Buf[61].Feature_n = FeatureBuf_747;
         Mult_Buf[61].Weight_n = Wgt_2_747;
         Mult_Buf[62].Feature_n = FeatureBuf_748;
         Mult_Buf[62].Weight_n = Wgt_2_748;
         Mult_Buf[63].Feature_n = FeatureBuf_749;
         Mult_Buf[63].Weight_n = Wgt_2_749;
         Mult_Buf[64].Feature_n = FeatureBuf_750;
         Mult_Buf[64].Weight_n = Wgt_2_750;
         Mult_Buf[65].Feature_n = FeatureBuf_751;
         Mult_Buf[65].Weight_n = Wgt_2_751;
         Mult_Buf[66].Feature_n = FeatureBuf_752;
         Mult_Buf[66].Weight_n = Wgt_2_752;
         Mult_Buf[67].Feature_n = FeatureBuf_753;
         Mult_Buf[67].Weight_n = Wgt_2_753;
         Mult_Buf[68].Feature_n = FeatureBuf_754;
         Mult_Buf[68].Weight_n = Wgt_2_754;
         Mult_Buf[69].Feature_n = FeatureBuf_755;
         Mult_Buf[69].Weight_n = Wgt_2_755;
         Mult_Buf[70].Feature_n = FeatureBuf_756;
         Mult_Buf[70].Weight_n = Wgt_2_756;
         Mult_Buf[71].Feature_n = FeatureBuf_757;
         Mult_Buf[71].Weight_n = Wgt_2_757;
         Mult_Buf[72].Feature_n = FeatureBuf_758;
         Mult_Buf[72].Weight_n = Wgt_2_758;
         Mult_Buf[73].Feature_n = FeatureBuf_759;
         Mult_Buf[73].Weight_n = Wgt_2_759;
         Mult_Buf[74].Feature_n = FeatureBuf_760;
         Mult_Buf[74].Weight_n = Wgt_2_760;
         Mult_Buf[75].Feature_n = FeatureBuf_761;
         Mult_Buf[75].Weight_n = Wgt_2_761;
         Mult_Buf[76].Feature_n = FeatureBuf_762;
         Mult_Buf[76].Weight_n = Wgt_2_762;
         Mult_Buf[77].Feature_n = FeatureBuf_763;
         Mult_Buf[77].Weight_n = Wgt_2_763;
         Mult_Buf[78].Feature_n = FeatureBuf_764;
         Mult_Buf[78].Weight_n = Wgt_2_764;
         Mult_Buf[79].Feature_n = FeatureBuf_765;
         Mult_Buf[79].Weight_n = Wgt_2_765;
         Mult_Buf[80].Feature_n = FeatureBuf_766;
         Mult_Buf[80].Weight_n = Wgt_2_766;
         Mult_Buf[81].Feature_n = FeatureBuf_767;
         Mult_Buf[81].Weight_n = Wgt_2_767;
         Mult_Buf[82].Feature_n = FeatureBuf_768;
         Mult_Buf[82].Weight_n = Wgt_2_768;
         Mult_Buf[83].Feature_n = FeatureBuf_769;
         Mult_Buf[83].Weight_n = Wgt_2_769;
         Mult_Buf[84].Feature_n = FeatureBuf_770;
         Mult_Buf[84].Weight_n = Wgt_2_770;
         Mult_Buf[85].Feature_n = FeatureBuf_771;
         Mult_Buf[85].Weight_n = Wgt_2_771;
         Mult_Buf[86].Feature_n = FeatureBuf_772;
         Mult_Buf[86].Weight_n = Wgt_2_772;
         Mult_Buf[87].Feature_n = FeatureBuf_773;
         Mult_Buf[87].Weight_n = Wgt_2_773;
         Mult_Buf[88].Feature_n = FeatureBuf_774;
         Mult_Buf[88].Weight_n = Wgt_2_774;
         Mult_Buf[89].Feature_n = FeatureBuf_775;
         Mult_Buf[89].Weight_n = Wgt_2_775;
         Mult_Buf[90].Feature_n = FeatureBuf_776;
         Mult_Buf[90].Weight_n = Wgt_2_776;
         Mult_Buf[91].Feature_n = FeatureBuf_777;
         Mult_Buf[91].Weight_n = Wgt_2_777;
         Mult_Buf[92].Feature_n = FeatureBuf_778;
         Mult_Buf[92].Weight_n = Wgt_2_778;
         Mult_Buf[93].Feature_n = FeatureBuf_779;
         Mult_Buf[93].Weight_n = Wgt_2_779;
         Mult_Buf[94].Feature_n = FeatureBuf_780;
         Mult_Buf[94].Weight_n = Wgt_2_780;
         Mult_Buf[95].Feature_n = FeatureBuf_781;
         Mult_Buf[95].Weight_n = Wgt_2_781;
         Mult_Buf[96].Feature_n = FeatureBuf_782;
         Mult_Buf[96].Weight_n = Wgt_2_782;
         Mult_Buf[97].Feature_n = FeatureBuf_783;
         Mult_Buf[97].Weight_n = Wgt_2_783;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     //Collect Partial result form Adder
         Res_0_1_n = Part_Res;
     end
    26:begin
     nxt_state = 27;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_0;
         Mult_Buf[0].Weight_n = Wgt_3_0;
         Mult_Buf[1].Feature_n = FeatureBuf_1;
         Mult_Buf[1].Weight_n = Wgt_3_1;
         Mult_Buf[2].Feature_n = FeatureBuf_2;
         Mult_Buf[2].Weight_n = Wgt_3_2;
         Mult_Buf[3].Feature_n = FeatureBuf_3;
         Mult_Buf[3].Weight_n = Wgt_3_3;
         Mult_Buf[4].Feature_n = FeatureBuf_4;
         Mult_Buf[4].Weight_n = Wgt_3_4;
         Mult_Buf[5].Feature_n = FeatureBuf_5;
         Mult_Buf[5].Weight_n = Wgt_3_5;
         Mult_Buf[6].Feature_n = FeatureBuf_6;
         Mult_Buf[6].Weight_n = Wgt_3_6;
         Mult_Buf[7].Feature_n = FeatureBuf_7;
         Mult_Buf[7].Weight_n = Wgt_3_7;
         Mult_Buf[8].Feature_n = FeatureBuf_8;
         Mult_Buf[8].Weight_n = Wgt_3_8;
         Mult_Buf[9].Feature_n = FeatureBuf_9;
         Mult_Buf[9].Weight_n = Wgt_3_9;
         Mult_Buf[10].Feature_n = FeatureBuf_10;
         Mult_Buf[10].Weight_n = Wgt_3_10;
         Mult_Buf[11].Feature_n = FeatureBuf_11;
         Mult_Buf[11].Weight_n = Wgt_3_11;
         Mult_Buf[12].Feature_n = FeatureBuf_12;
         Mult_Buf[12].Weight_n = Wgt_3_12;
         Mult_Buf[13].Feature_n = FeatureBuf_13;
         Mult_Buf[13].Weight_n = Wgt_3_13;
         Mult_Buf[14].Feature_n = FeatureBuf_14;
         Mult_Buf[14].Weight_n = Wgt_3_14;
         Mult_Buf[15].Feature_n = FeatureBuf_15;
         Mult_Buf[15].Weight_n = Wgt_3_15;
         Mult_Buf[16].Feature_n = FeatureBuf_16;
         Mult_Buf[16].Weight_n = Wgt_3_16;
         Mult_Buf[17].Feature_n = FeatureBuf_17;
         Mult_Buf[17].Weight_n = Wgt_3_17;
         Mult_Buf[18].Feature_n = FeatureBuf_18;
         Mult_Buf[18].Weight_n = Wgt_3_18;
         Mult_Buf[19].Feature_n = FeatureBuf_19;
         Mult_Buf[19].Weight_n = Wgt_3_19;
         Mult_Buf[20].Feature_n = FeatureBuf_20;
         Mult_Buf[20].Weight_n = Wgt_3_20;
         Mult_Buf[21].Feature_n = FeatureBuf_21;
         Mult_Buf[21].Weight_n = Wgt_3_21;
         Mult_Buf[22].Feature_n = FeatureBuf_22;
         Mult_Buf[22].Weight_n = Wgt_3_22;
         Mult_Buf[23].Feature_n = FeatureBuf_23;
         Mult_Buf[23].Weight_n = Wgt_3_23;
         Mult_Buf[24].Feature_n = FeatureBuf_24;
         Mult_Buf[24].Weight_n = Wgt_3_24;
         Mult_Buf[25].Feature_n = FeatureBuf_25;
         Mult_Buf[25].Weight_n = Wgt_3_25;
         Mult_Buf[26].Feature_n = FeatureBuf_26;
         Mult_Buf[26].Weight_n = Wgt_3_26;
         Mult_Buf[27].Feature_n = FeatureBuf_27;
         Mult_Buf[27].Weight_n = Wgt_3_27;
         Mult_Buf[28].Feature_n = FeatureBuf_28;
         Mult_Buf[28].Weight_n = Wgt_3_28;
         Mult_Buf[29].Feature_n = FeatureBuf_29;
         Mult_Buf[29].Weight_n = Wgt_3_29;
         Mult_Buf[30].Feature_n = FeatureBuf_30;
         Mult_Buf[30].Weight_n = Wgt_3_30;
         Mult_Buf[31].Feature_n = FeatureBuf_31;
         Mult_Buf[31].Weight_n = Wgt_3_31;
         Mult_Buf[32].Feature_n = FeatureBuf_32;
         Mult_Buf[32].Weight_n = Wgt_3_32;
         Mult_Buf[33].Feature_n = FeatureBuf_33;
         Mult_Buf[33].Weight_n = Wgt_3_33;
         Mult_Buf[34].Feature_n = FeatureBuf_34;
         Mult_Buf[34].Weight_n = Wgt_3_34;
         Mult_Buf[35].Feature_n = FeatureBuf_35;
         Mult_Buf[35].Weight_n = Wgt_3_35;
         Mult_Buf[36].Feature_n = FeatureBuf_36;
         Mult_Buf[36].Weight_n = Wgt_3_36;
         Mult_Buf[37].Feature_n = FeatureBuf_37;
         Mult_Buf[37].Weight_n = Wgt_3_37;
         Mult_Buf[38].Feature_n = FeatureBuf_38;
         Mult_Buf[38].Weight_n = Wgt_3_38;
         Mult_Buf[39].Feature_n = FeatureBuf_39;
         Mult_Buf[39].Weight_n = Wgt_3_39;
         Mult_Buf[40].Feature_n = FeatureBuf_40;
         Mult_Buf[40].Weight_n = Wgt_3_40;
         Mult_Buf[41].Feature_n = FeatureBuf_41;
         Mult_Buf[41].Weight_n = Wgt_3_41;
         Mult_Buf[42].Feature_n = FeatureBuf_42;
         Mult_Buf[42].Weight_n = Wgt_3_42;
         Mult_Buf[43].Feature_n = FeatureBuf_43;
         Mult_Buf[43].Weight_n = Wgt_3_43;
         Mult_Buf[44].Feature_n = FeatureBuf_44;
         Mult_Buf[44].Weight_n = Wgt_3_44;
         Mult_Buf[45].Feature_n = FeatureBuf_45;
         Mult_Buf[45].Weight_n = Wgt_3_45;
         Mult_Buf[46].Feature_n = FeatureBuf_46;
         Mult_Buf[46].Weight_n = Wgt_3_46;
         Mult_Buf[47].Feature_n = FeatureBuf_47;
         Mult_Buf[47].Weight_n = Wgt_3_47;
         Mult_Buf[48].Feature_n = FeatureBuf_48;
         Mult_Buf[48].Weight_n = Wgt_3_48;
         Mult_Buf[49].Feature_n = FeatureBuf_49;
         Mult_Buf[49].Weight_n = Wgt_3_49;
         Mult_Buf[50].Feature_n = FeatureBuf_50;
         Mult_Buf[50].Weight_n = Wgt_3_50;
         Mult_Buf[51].Feature_n = FeatureBuf_51;
         Mult_Buf[51].Weight_n = Wgt_3_51;
         Mult_Buf[52].Feature_n = FeatureBuf_52;
         Mult_Buf[52].Weight_n = Wgt_3_52;
         Mult_Buf[53].Feature_n = FeatureBuf_53;
         Mult_Buf[53].Weight_n = Wgt_3_53;
         Mult_Buf[54].Feature_n = FeatureBuf_54;
         Mult_Buf[54].Weight_n = Wgt_3_54;
         Mult_Buf[55].Feature_n = FeatureBuf_55;
         Mult_Buf[55].Weight_n = Wgt_3_55;
         Mult_Buf[56].Feature_n = FeatureBuf_56;
         Mult_Buf[56].Weight_n = Wgt_3_56;
         Mult_Buf[57].Feature_n = FeatureBuf_57;
         Mult_Buf[57].Weight_n = Wgt_3_57;
         Mult_Buf[58].Feature_n = FeatureBuf_58;
         Mult_Buf[58].Weight_n = Wgt_3_58;
         Mult_Buf[59].Feature_n = FeatureBuf_59;
         Mult_Buf[59].Weight_n = Wgt_3_59;
         Mult_Buf[60].Feature_n = FeatureBuf_60;
         Mult_Buf[60].Weight_n = Wgt_3_60;
         Mult_Buf[61].Feature_n = FeatureBuf_61;
         Mult_Buf[61].Weight_n = Wgt_3_61;
         Mult_Buf[62].Feature_n = FeatureBuf_62;
         Mult_Buf[62].Weight_n = Wgt_3_62;
         Mult_Buf[63].Feature_n = FeatureBuf_63;
         Mult_Buf[63].Weight_n = Wgt_3_63;
         Mult_Buf[64].Feature_n = FeatureBuf_64;
         Mult_Buf[64].Weight_n = Wgt_3_64;
         Mult_Buf[65].Feature_n = FeatureBuf_65;
         Mult_Buf[65].Weight_n = Wgt_3_65;
         Mult_Buf[66].Feature_n = FeatureBuf_66;
         Mult_Buf[66].Weight_n = Wgt_3_66;
         Mult_Buf[67].Feature_n = FeatureBuf_67;
         Mult_Buf[67].Weight_n = Wgt_3_67;
         Mult_Buf[68].Feature_n = FeatureBuf_68;
         Mult_Buf[68].Weight_n = Wgt_3_68;
         Mult_Buf[69].Feature_n = FeatureBuf_69;
         Mult_Buf[69].Weight_n = Wgt_3_69;
         Mult_Buf[70].Feature_n = FeatureBuf_70;
         Mult_Buf[70].Weight_n = Wgt_3_70;
         Mult_Buf[71].Feature_n = FeatureBuf_71;
         Mult_Buf[71].Weight_n = Wgt_3_71;
         Mult_Buf[72].Feature_n = FeatureBuf_72;
         Mult_Buf[72].Weight_n = Wgt_3_72;
         Mult_Buf[73].Feature_n = FeatureBuf_73;
         Mult_Buf[73].Weight_n = Wgt_3_73;
         Mult_Buf[74].Feature_n = FeatureBuf_74;
         Mult_Buf[74].Weight_n = Wgt_3_74;
         Mult_Buf[75].Feature_n = FeatureBuf_75;
         Mult_Buf[75].Weight_n = Wgt_3_75;
         Mult_Buf[76].Feature_n = FeatureBuf_76;
         Mult_Buf[76].Weight_n = Wgt_3_76;
         Mult_Buf[77].Feature_n = FeatureBuf_77;
         Mult_Buf[77].Weight_n = Wgt_3_77;
         Mult_Buf[78].Feature_n = FeatureBuf_78;
         Mult_Buf[78].Weight_n = Wgt_3_78;
         Mult_Buf[79].Feature_n = FeatureBuf_79;
         Mult_Buf[79].Weight_n = Wgt_3_79;
         Mult_Buf[80].Feature_n = FeatureBuf_80;
         Mult_Buf[80].Weight_n = Wgt_3_80;
         Mult_Buf[81].Feature_n = FeatureBuf_81;
         Mult_Buf[81].Weight_n = Wgt_3_81;
         Mult_Buf[82].Feature_n = FeatureBuf_82;
         Mult_Buf[82].Weight_n = Wgt_3_82;
         Mult_Buf[83].Feature_n = FeatureBuf_83;
         Mult_Buf[83].Weight_n = Wgt_3_83;
         Mult_Buf[84].Feature_n = FeatureBuf_84;
         Mult_Buf[84].Weight_n = Wgt_3_84;
         Mult_Buf[85].Feature_n = FeatureBuf_85;
         Mult_Buf[85].Weight_n = Wgt_3_85;
         Mult_Buf[86].Feature_n = FeatureBuf_86;
         Mult_Buf[86].Weight_n = Wgt_3_86;
         Mult_Buf[87].Feature_n = FeatureBuf_87;
         Mult_Buf[87].Weight_n = Wgt_3_87;
         Mult_Buf[88].Feature_n = FeatureBuf_88;
         Mult_Buf[88].Weight_n = Wgt_3_88;
         Mult_Buf[89].Feature_n = FeatureBuf_89;
         Mult_Buf[89].Weight_n = Wgt_3_89;
         Mult_Buf[90].Feature_n = FeatureBuf_90;
         Mult_Buf[90].Weight_n = Wgt_3_90;
         Mult_Buf[91].Feature_n = FeatureBuf_91;
         Mult_Buf[91].Weight_n = Wgt_3_91;
         Mult_Buf[92].Feature_n = FeatureBuf_92;
         Mult_Buf[92].Weight_n = Wgt_3_92;
         Mult_Buf[93].Feature_n = FeatureBuf_93;
         Mult_Buf[93].Weight_n = Wgt_3_93;
         Mult_Buf[94].Feature_n = FeatureBuf_94;
         Mult_Buf[94].Weight_n = Wgt_3_94;
         Mult_Buf[95].Feature_n = FeatureBuf_95;
         Mult_Buf[95].Weight_n = Wgt_3_95;
         Mult_Buf[96].Feature_n = FeatureBuf_96;
         Mult_Buf[96].Weight_n = Wgt_3_96;
         Mult_Buf[97].Feature_n = FeatureBuf_97;
         Mult_Buf[97].Weight_n = Wgt_3_97;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     //Collect Partial result form Adder
         Res_0_2_n = Part_Res;
     end
    27:begin
     nxt_state = 28;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_98;
         Mult_Buf[0].Weight_n = Wgt_3_98;
         Mult_Buf[1].Feature_n = FeatureBuf_99;
         Mult_Buf[1].Weight_n = Wgt_3_99;
         Mult_Buf[2].Feature_n = FeatureBuf_100;
         Mult_Buf[2].Weight_n = Wgt_3_100;
         Mult_Buf[3].Feature_n = FeatureBuf_101;
         Mult_Buf[3].Weight_n = Wgt_3_101;
         Mult_Buf[4].Feature_n = FeatureBuf_102;
         Mult_Buf[4].Weight_n = Wgt_3_102;
         Mult_Buf[5].Feature_n = FeatureBuf_103;
         Mult_Buf[5].Weight_n = Wgt_3_103;
         Mult_Buf[6].Feature_n = FeatureBuf_104;
         Mult_Buf[6].Weight_n = Wgt_3_104;
         Mult_Buf[7].Feature_n = FeatureBuf_105;
         Mult_Buf[7].Weight_n = Wgt_3_105;
         Mult_Buf[8].Feature_n = FeatureBuf_106;
         Mult_Buf[8].Weight_n = Wgt_3_106;
         Mult_Buf[9].Feature_n = FeatureBuf_107;
         Mult_Buf[9].Weight_n = Wgt_3_107;
         Mult_Buf[10].Feature_n = FeatureBuf_108;
         Mult_Buf[10].Weight_n = Wgt_3_108;
         Mult_Buf[11].Feature_n = FeatureBuf_109;
         Mult_Buf[11].Weight_n = Wgt_3_109;
         Mult_Buf[12].Feature_n = FeatureBuf_110;
         Mult_Buf[12].Weight_n = Wgt_3_110;
         Mult_Buf[13].Feature_n = FeatureBuf_111;
         Mult_Buf[13].Weight_n = Wgt_3_111;
         Mult_Buf[14].Feature_n = FeatureBuf_112;
         Mult_Buf[14].Weight_n = Wgt_3_112;
         Mult_Buf[15].Feature_n = FeatureBuf_113;
         Mult_Buf[15].Weight_n = Wgt_3_113;
         Mult_Buf[16].Feature_n = FeatureBuf_114;
         Mult_Buf[16].Weight_n = Wgt_3_114;
         Mult_Buf[17].Feature_n = FeatureBuf_115;
         Mult_Buf[17].Weight_n = Wgt_3_115;
         Mult_Buf[18].Feature_n = FeatureBuf_116;
         Mult_Buf[18].Weight_n = Wgt_3_116;
         Mult_Buf[19].Feature_n = FeatureBuf_117;
         Mult_Buf[19].Weight_n = Wgt_3_117;
         Mult_Buf[20].Feature_n = FeatureBuf_118;
         Mult_Buf[20].Weight_n = Wgt_3_118;
         Mult_Buf[21].Feature_n = FeatureBuf_119;
         Mult_Buf[21].Weight_n = Wgt_3_119;
         Mult_Buf[22].Feature_n = FeatureBuf_120;
         Mult_Buf[22].Weight_n = Wgt_3_120;
         Mult_Buf[23].Feature_n = FeatureBuf_121;
         Mult_Buf[23].Weight_n = Wgt_3_121;
         Mult_Buf[24].Feature_n = FeatureBuf_122;
         Mult_Buf[24].Weight_n = Wgt_3_122;
         Mult_Buf[25].Feature_n = FeatureBuf_123;
         Mult_Buf[25].Weight_n = Wgt_3_123;
         Mult_Buf[26].Feature_n = FeatureBuf_124;
         Mult_Buf[26].Weight_n = Wgt_3_124;
         Mult_Buf[27].Feature_n = FeatureBuf_125;
         Mult_Buf[27].Weight_n = Wgt_3_125;
         Mult_Buf[28].Feature_n = FeatureBuf_126;
         Mult_Buf[28].Weight_n = Wgt_3_126;
         Mult_Buf[29].Feature_n = FeatureBuf_127;
         Mult_Buf[29].Weight_n = Wgt_3_127;
         Mult_Buf[30].Feature_n = FeatureBuf_128;
         Mult_Buf[30].Weight_n = Wgt_3_128;
         Mult_Buf[31].Feature_n = FeatureBuf_129;
         Mult_Buf[31].Weight_n = Wgt_3_129;
         Mult_Buf[32].Feature_n = FeatureBuf_130;
         Mult_Buf[32].Weight_n = Wgt_3_130;
         Mult_Buf[33].Feature_n = FeatureBuf_131;
         Mult_Buf[33].Weight_n = Wgt_3_131;
         Mult_Buf[34].Feature_n = FeatureBuf_132;
         Mult_Buf[34].Weight_n = Wgt_3_132;
         Mult_Buf[35].Feature_n = FeatureBuf_133;
         Mult_Buf[35].Weight_n = Wgt_3_133;
         Mult_Buf[36].Feature_n = FeatureBuf_134;
         Mult_Buf[36].Weight_n = Wgt_3_134;
         Mult_Buf[37].Feature_n = FeatureBuf_135;
         Mult_Buf[37].Weight_n = Wgt_3_135;
         Mult_Buf[38].Feature_n = FeatureBuf_136;
         Mult_Buf[38].Weight_n = Wgt_3_136;
         Mult_Buf[39].Feature_n = FeatureBuf_137;
         Mult_Buf[39].Weight_n = Wgt_3_137;
         Mult_Buf[40].Feature_n = FeatureBuf_138;
         Mult_Buf[40].Weight_n = Wgt_3_138;
         Mult_Buf[41].Feature_n = FeatureBuf_139;
         Mult_Buf[41].Weight_n = Wgt_3_139;
         Mult_Buf[42].Feature_n = FeatureBuf_140;
         Mult_Buf[42].Weight_n = Wgt_3_140;
         Mult_Buf[43].Feature_n = FeatureBuf_141;
         Mult_Buf[43].Weight_n = Wgt_3_141;
         Mult_Buf[44].Feature_n = FeatureBuf_142;
         Mult_Buf[44].Weight_n = Wgt_3_142;
         Mult_Buf[45].Feature_n = FeatureBuf_143;
         Mult_Buf[45].Weight_n = Wgt_3_143;
         Mult_Buf[46].Feature_n = FeatureBuf_144;
         Mult_Buf[46].Weight_n = Wgt_3_144;
         Mult_Buf[47].Feature_n = FeatureBuf_145;
         Mult_Buf[47].Weight_n = Wgt_3_145;
         Mult_Buf[48].Feature_n = FeatureBuf_146;
         Mult_Buf[48].Weight_n = Wgt_3_146;
         Mult_Buf[49].Feature_n = FeatureBuf_147;
         Mult_Buf[49].Weight_n = Wgt_3_147;
         Mult_Buf[50].Feature_n = FeatureBuf_148;
         Mult_Buf[50].Weight_n = Wgt_3_148;
         Mult_Buf[51].Feature_n = FeatureBuf_149;
         Mult_Buf[51].Weight_n = Wgt_3_149;
         Mult_Buf[52].Feature_n = FeatureBuf_150;
         Mult_Buf[52].Weight_n = Wgt_3_150;
         Mult_Buf[53].Feature_n = FeatureBuf_151;
         Mult_Buf[53].Weight_n = Wgt_3_151;
         Mult_Buf[54].Feature_n = FeatureBuf_152;
         Mult_Buf[54].Weight_n = Wgt_3_152;
         Mult_Buf[55].Feature_n = FeatureBuf_153;
         Mult_Buf[55].Weight_n = Wgt_3_153;
         Mult_Buf[56].Feature_n = FeatureBuf_154;
         Mult_Buf[56].Weight_n = Wgt_3_154;
         Mult_Buf[57].Feature_n = FeatureBuf_155;
         Mult_Buf[57].Weight_n = Wgt_3_155;
         Mult_Buf[58].Feature_n = FeatureBuf_156;
         Mult_Buf[58].Weight_n = Wgt_3_156;
         Mult_Buf[59].Feature_n = FeatureBuf_157;
         Mult_Buf[59].Weight_n = Wgt_3_157;
         Mult_Buf[60].Feature_n = FeatureBuf_158;
         Mult_Buf[60].Weight_n = Wgt_3_158;
         Mult_Buf[61].Feature_n = FeatureBuf_159;
         Mult_Buf[61].Weight_n = Wgt_3_159;
         Mult_Buf[62].Feature_n = FeatureBuf_160;
         Mult_Buf[62].Weight_n = Wgt_3_160;
         Mult_Buf[63].Feature_n = FeatureBuf_161;
         Mult_Buf[63].Weight_n = Wgt_3_161;
         Mult_Buf[64].Feature_n = FeatureBuf_162;
         Mult_Buf[64].Weight_n = Wgt_3_162;
         Mult_Buf[65].Feature_n = FeatureBuf_163;
         Mult_Buf[65].Weight_n = Wgt_3_163;
         Mult_Buf[66].Feature_n = FeatureBuf_164;
         Mult_Buf[66].Weight_n = Wgt_3_164;
         Mult_Buf[67].Feature_n = FeatureBuf_165;
         Mult_Buf[67].Weight_n = Wgt_3_165;
         Mult_Buf[68].Feature_n = FeatureBuf_166;
         Mult_Buf[68].Weight_n = Wgt_3_166;
         Mult_Buf[69].Feature_n = FeatureBuf_167;
         Mult_Buf[69].Weight_n = Wgt_3_167;
         Mult_Buf[70].Feature_n = FeatureBuf_168;
         Mult_Buf[70].Weight_n = Wgt_3_168;
         Mult_Buf[71].Feature_n = FeatureBuf_169;
         Mult_Buf[71].Weight_n = Wgt_3_169;
         Mult_Buf[72].Feature_n = FeatureBuf_170;
         Mult_Buf[72].Weight_n = Wgt_3_170;
         Mult_Buf[73].Feature_n = FeatureBuf_171;
         Mult_Buf[73].Weight_n = Wgt_3_171;
         Mult_Buf[74].Feature_n = FeatureBuf_172;
         Mult_Buf[74].Weight_n = Wgt_3_172;
         Mult_Buf[75].Feature_n = FeatureBuf_173;
         Mult_Buf[75].Weight_n = Wgt_3_173;
         Mult_Buf[76].Feature_n = FeatureBuf_174;
         Mult_Buf[76].Weight_n = Wgt_3_174;
         Mult_Buf[77].Feature_n = FeatureBuf_175;
         Mult_Buf[77].Weight_n = Wgt_3_175;
         Mult_Buf[78].Feature_n = FeatureBuf_176;
         Mult_Buf[78].Weight_n = Wgt_3_176;
         Mult_Buf[79].Feature_n = FeatureBuf_177;
         Mult_Buf[79].Weight_n = Wgt_3_177;
         Mult_Buf[80].Feature_n = FeatureBuf_178;
         Mult_Buf[80].Weight_n = Wgt_3_178;
         Mult_Buf[81].Feature_n = FeatureBuf_179;
         Mult_Buf[81].Weight_n = Wgt_3_179;
         Mult_Buf[82].Feature_n = FeatureBuf_180;
         Mult_Buf[82].Weight_n = Wgt_3_180;
         Mult_Buf[83].Feature_n = FeatureBuf_181;
         Mult_Buf[83].Weight_n = Wgt_3_181;
         Mult_Buf[84].Feature_n = FeatureBuf_182;
         Mult_Buf[84].Weight_n = Wgt_3_182;
         Mult_Buf[85].Feature_n = FeatureBuf_183;
         Mult_Buf[85].Weight_n = Wgt_3_183;
         Mult_Buf[86].Feature_n = FeatureBuf_184;
         Mult_Buf[86].Weight_n = Wgt_3_184;
         Mult_Buf[87].Feature_n = FeatureBuf_185;
         Mult_Buf[87].Weight_n = Wgt_3_185;
         Mult_Buf[88].Feature_n = FeatureBuf_186;
         Mult_Buf[88].Weight_n = Wgt_3_186;
         Mult_Buf[89].Feature_n = FeatureBuf_187;
         Mult_Buf[89].Weight_n = Wgt_3_187;
         Mult_Buf[90].Feature_n = FeatureBuf_188;
         Mult_Buf[90].Weight_n = Wgt_3_188;
         Mult_Buf[91].Feature_n = FeatureBuf_189;
         Mult_Buf[91].Weight_n = Wgt_3_189;
         Mult_Buf[92].Feature_n = FeatureBuf_190;
         Mult_Buf[92].Weight_n = Wgt_3_190;
         Mult_Buf[93].Feature_n = FeatureBuf_191;
         Mult_Buf[93].Weight_n = Wgt_3_191;
         Mult_Buf[94].Feature_n = FeatureBuf_192;
         Mult_Buf[94].Weight_n = Wgt_3_192;
         Mult_Buf[95].Feature_n = FeatureBuf_193;
         Mult_Buf[95].Weight_n = Wgt_3_193;
         Mult_Buf[96].Feature_n = FeatureBuf_194;
         Mult_Buf[96].Weight_n = Wgt_3_194;
         Mult_Buf[97].Feature_n = FeatureBuf_195;
         Mult_Buf[97].Weight_n = Wgt_3_195;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     //Collect Partial result form Adder
         Res_0_3_n = Part_Res;
     end
    28:begin
     nxt_state = 29;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_196;
         Mult_Buf[0].Weight_n = Wgt_3_196;
         Mult_Buf[1].Feature_n = FeatureBuf_197;
         Mult_Buf[1].Weight_n = Wgt_3_197;
         Mult_Buf[2].Feature_n = FeatureBuf_198;
         Mult_Buf[2].Weight_n = Wgt_3_198;
         Mult_Buf[3].Feature_n = FeatureBuf_199;
         Mult_Buf[3].Weight_n = Wgt_3_199;
         Mult_Buf[4].Feature_n = FeatureBuf_200;
         Mult_Buf[4].Weight_n = Wgt_3_200;
         Mult_Buf[5].Feature_n = FeatureBuf_201;
         Mult_Buf[5].Weight_n = Wgt_3_201;
         Mult_Buf[6].Feature_n = FeatureBuf_202;
         Mult_Buf[6].Weight_n = Wgt_3_202;
         Mult_Buf[7].Feature_n = FeatureBuf_203;
         Mult_Buf[7].Weight_n = Wgt_3_203;
         Mult_Buf[8].Feature_n = FeatureBuf_204;
         Mult_Buf[8].Weight_n = Wgt_3_204;
         Mult_Buf[9].Feature_n = FeatureBuf_205;
         Mult_Buf[9].Weight_n = Wgt_3_205;
         Mult_Buf[10].Feature_n = FeatureBuf_206;
         Mult_Buf[10].Weight_n = Wgt_3_206;
         Mult_Buf[11].Feature_n = FeatureBuf_207;
         Mult_Buf[11].Weight_n = Wgt_3_207;
         Mult_Buf[12].Feature_n = FeatureBuf_208;
         Mult_Buf[12].Weight_n = Wgt_3_208;
         Mult_Buf[13].Feature_n = FeatureBuf_209;
         Mult_Buf[13].Weight_n = Wgt_3_209;
         Mult_Buf[14].Feature_n = FeatureBuf_210;
         Mult_Buf[14].Weight_n = Wgt_3_210;
         Mult_Buf[15].Feature_n = FeatureBuf_211;
         Mult_Buf[15].Weight_n = Wgt_3_211;
         Mult_Buf[16].Feature_n = FeatureBuf_212;
         Mult_Buf[16].Weight_n = Wgt_3_212;
         Mult_Buf[17].Feature_n = FeatureBuf_213;
         Mult_Buf[17].Weight_n = Wgt_3_213;
         Mult_Buf[18].Feature_n = FeatureBuf_214;
         Mult_Buf[18].Weight_n = Wgt_3_214;
         Mult_Buf[19].Feature_n = FeatureBuf_215;
         Mult_Buf[19].Weight_n = Wgt_3_215;
         Mult_Buf[20].Feature_n = FeatureBuf_216;
         Mult_Buf[20].Weight_n = Wgt_3_216;
         Mult_Buf[21].Feature_n = FeatureBuf_217;
         Mult_Buf[21].Weight_n = Wgt_3_217;
         Mult_Buf[22].Feature_n = FeatureBuf_218;
         Mult_Buf[22].Weight_n = Wgt_3_218;
         Mult_Buf[23].Feature_n = FeatureBuf_219;
         Mult_Buf[23].Weight_n = Wgt_3_219;
         Mult_Buf[24].Feature_n = FeatureBuf_220;
         Mult_Buf[24].Weight_n = Wgt_3_220;
         Mult_Buf[25].Feature_n = FeatureBuf_221;
         Mult_Buf[25].Weight_n = Wgt_3_221;
         Mult_Buf[26].Feature_n = FeatureBuf_222;
         Mult_Buf[26].Weight_n = Wgt_3_222;
         Mult_Buf[27].Feature_n = FeatureBuf_223;
         Mult_Buf[27].Weight_n = Wgt_3_223;
         Mult_Buf[28].Feature_n = FeatureBuf_224;
         Mult_Buf[28].Weight_n = Wgt_3_224;
         Mult_Buf[29].Feature_n = FeatureBuf_225;
         Mult_Buf[29].Weight_n = Wgt_3_225;
         Mult_Buf[30].Feature_n = FeatureBuf_226;
         Mult_Buf[30].Weight_n = Wgt_3_226;
         Mult_Buf[31].Feature_n = FeatureBuf_227;
         Mult_Buf[31].Weight_n = Wgt_3_227;
         Mult_Buf[32].Feature_n = FeatureBuf_228;
         Mult_Buf[32].Weight_n = Wgt_3_228;
         Mult_Buf[33].Feature_n = FeatureBuf_229;
         Mult_Buf[33].Weight_n = Wgt_3_229;
         Mult_Buf[34].Feature_n = FeatureBuf_230;
         Mult_Buf[34].Weight_n = Wgt_3_230;
         Mult_Buf[35].Feature_n = FeatureBuf_231;
         Mult_Buf[35].Weight_n = Wgt_3_231;
         Mult_Buf[36].Feature_n = FeatureBuf_232;
         Mult_Buf[36].Weight_n = Wgt_3_232;
         Mult_Buf[37].Feature_n = FeatureBuf_233;
         Mult_Buf[37].Weight_n = Wgt_3_233;
         Mult_Buf[38].Feature_n = FeatureBuf_234;
         Mult_Buf[38].Weight_n = Wgt_3_234;
         Mult_Buf[39].Feature_n = FeatureBuf_235;
         Mult_Buf[39].Weight_n = Wgt_3_235;
         Mult_Buf[40].Feature_n = FeatureBuf_236;
         Mult_Buf[40].Weight_n = Wgt_3_236;
         Mult_Buf[41].Feature_n = FeatureBuf_237;
         Mult_Buf[41].Weight_n = Wgt_3_237;
         Mult_Buf[42].Feature_n = FeatureBuf_238;
         Mult_Buf[42].Weight_n = Wgt_3_238;
         Mult_Buf[43].Feature_n = FeatureBuf_239;
         Mult_Buf[43].Weight_n = Wgt_3_239;
         Mult_Buf[44].Feature_n = FeatureBuf_240;
         Mult_Buf[44].Weight_n = Wgt_3_240;
         Mult_Buf[45].Feature_n = FeatureBuf_241;
         Mult_Buf[45].Weight_n = Wgt_3_241;
         Mult_Buf[46].Feature_n = FeatureBuf_242;
         Mult_Buf[46].Weight_n = Wgt_3_242;
         Mult_Buf[47].Feature_n = FeatureBuf_243;
         Mult_Buf[47].Weight_n = Wgt_3_243;
         Mult_Buf[48].Feature_n = FeatureBuf_244;
         Mult_Buf[48].Weight_n = Wgt_3_244;
         Mult_Buf[49].Feature_n = FeatureBuf_245;
         Mult_Buf[49].Weight_n = Wgt_3_245;
         Mult_Buf[50].Feature_n = FeatureBuf_246;
         Mult_Buf[50].Weight_n = Wgt_3_246;
         Mult_Buf[51].Feature_n = FeatureBuf_247;
         Mult_Buf[51].Weight_n = Wgt_3_247;
         Mult_Buf[52].Feature_n = FeatureBuf_248;
         Mult_Buf[52].Weight_n = Wgt_3_248;
         Mult_Buf[53].Feature_n = FeatureBuf_249;
         Mult_Buf[53].Weight_n = Wgt_3_249;
         Mult_Buf[54].Feature_n = FeatureBuf_250;
         Mult_Buf[54].Weight_n = Wgt_3_250;
         Mult_Buf[55].Feature_n = FeatureBuf_251;
         Mult_Buf[55].Weight_n = Wgt_3_251;
         Mult_Buf[56].Feature_n = FeatureBuf_252;
         Mult_Buf[56].Weight_n = Wgt_3_252;
         Mult_Buf[57].Feature_n = FeatureBuf_253;
         Mult_Buf[57].Weight_n = Wgt_3_253;
         Mult_Buf[58].Feature_n = FeatureBuf_254;
         Mult_Buf[58].Weight_n = Wgt_3_254;
         Mult_Buf[59].Feature_n = FeatureBuf_255;
         Mult_Buf[59].Weight_n = Wgt_3_255;
         Mult_Buf[60].Feature_n = FeatureBuf_256;
         Mult_Buf[60].Weight_n = Wgt_3_256;
         Mult_Buf[61].Feature_n = FeatureBuf_257;
         Mult_Buf[61].Weight_n = Wgt_3_257;
         Mult_Buf[62].Feature_n = FeatureBuf_258;
         Mult_Buf[62].Weight_n = Wgt_3_258;
         Mult_Buf[63].Feature_n = FeatureBuf_259;
         Mult_Buf[63].Weight_n = Wgt_3_259;
         Mult_Buf[64].Feature_n = FeatureBuf_260;
         Mult_Buf[64].Weight_n = Wgt_3_260;
         Mult_Buf[65].Feature_n = FeatureBuf_261;
         Mult_Buf[65].Weight_n = Wgt_3_261;
         Mult_Buf[66].Feature_n = FeatureBuf_262;
         Mult_Buf[66].Weight_n = Wgt_3_262;
         Mult_Buf[67].Feature_n = FeatureBuf_263;
         Mult_Buf[67].Weight_n = Wgt_3_263;
         Mult_Buf[68].Feature_n = FeatureBuf_264;
         Mult_Buf[68].Weight_n = Wgt_3_264;
         Mult_Buf[69].Feature_n = FeatureBuf_265;
         Mult_Buf[69].Weight_n = Wgt_3_265;
         Mult_Buf[70].Feature_n = FeatureBuf_266;
         Mult_Buf[70].Weight_n = Wgt_3_266;
         Mult_Buf[71].Feature_n = FeatureBuf_267;
         Mult_Buf[71].Weight_n = Wgt_3_267;
         Mult_Buf[72].Feature_n = FeatureBuf_268;
         Mult_Buf[72].Weight_n = Wgt_3_268;
         Mult_Buf[73].Feature_n = FeatureBuf_269;
         Mult_Buf[73].Weight_n = Wgt_3_269;
         Mult_Buf[74].Feature_n = FeatureBuf_270;
         Mult_Buf[74].Weight_n = Wgt_3_270;
         Mult_Buf[75].Feature_n = FeatureBuf_271;
         Mult_Buf[75].Weight_n = Wgt_3_271;
         Mult_Buf[76].Feature_n = FeatureBuf_272;
         Mult_Buf[76].Weight_n = Wgt_3_272;
         Mult_Buf[77].Feature_n = FeatureBuf_273;
         Mult_Buf[77].Weight_n = Wgt_3_273;
         Mult_Buf[78].Feature_n = FeatureBuf_274;
         Mult_Buf[78].Weight_n = Wgt_3_274;
         Mult_Buf[79].Feature_n = FeatureBuf_275;
         Mult_Buf[79].Weight_n = Wgt_3_275;
         Mult_Buf[80].Feature_n = FeatureBuf_276;
         Mult_Buf[80].Weight_n = Wgt_3_276;
         Mult_Buf[81].Feature_n = FeatureBuf_277;
         Mult_Buf[81].Weight_n = Wgt_3_277;
         Mult_Buf[82].Feature_n = FeatureBuf_278;
         Mult_Buf[82].Weight_n = Wgt_3_278;
         Mult_Buf[83].Feature_n = FeatureBuf_279;
         Mult_Buf[83].Weight_n = Wgt_3_279;
         Mult_Buf[84].Feature_n = FeatureBuf_280;
         Mult_Buf[84].Weight_n = Wgt_3_280;
         Mult_Buf[85].Feature_n = FeatureBuf_281;
         Mult_Buf[85].Weight_n = Wgt_3_281;
         Mult_Buf[86].Feature_n = FeatureBuf_282;
         Mult_Buf[86].Weight_n = Wgt_3_282;
         Mult_Buf[87].Feature_n = FeatureBuf_283;
         Mult_Buf[87].Weight_n = Wgt_3_283;
         Mult_Buf[88].Feature_n = FeatureBuf_284;
         Mult_Buf[88].Weight_n = Wgt_3_284;
         Mult_Buf[89].Feature_n = FeatureBuf_285;
         Mult_Buf[89].Weight_n = Wgt_3_285;
         Mult_Buf[90].Feature_n = FeatureBuf_286;
         Mult_Buf[90].Weight_n = Wgt_3_286;
         Mult_Buf[91].Feature_n = FeatureBuf_287;
         Mult_Buf[91].Weight_n = Wgt_3_287;
         Mult_Buf[92].Feature_n = FeatureBuf_288;
         Mult_Buf[92].Weight_n = Wgt_3_288;
         Mult_Buf[93].Feature_n = FeatureBuf_289;
         Mult_Buf[93].Weight_n = Wgt_3_289;
         Mult_Buf[94].Feature_n = FeatureBuf_290;
         Mult_Buf[94].Weight_n = Wgt_3_290;
         Mult_Buf[95].Feature_n = FeatureBuf_291;
         Mult_Buf[95].Weight_n = Wgt_3_291;
         Mult_Buf[96].Feature_n = FeatureBuf_292;
         Mult_Buf[96].Weight_n = Wgt_3_292;
         Mult_Buf[97].Feature_n = FeatureBuf_293;
         Mult_Buf[97].Weight_n = Wgt_3_293;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     //Collect Partial result form Adder
         Res_0_4_n = Part_Res;
     end
    29:begin
     nxt_state = 30;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_294;
         Mult_Buf[0].Weight_n = Wgt_3_294;
         Mult_Buf[1].Feature_n = FeatureBuf_295;
         Mult_Buf[1].Weight_n = Wgt_3_295;
         Mult_Buf[2].Feature_n = FeatureBuf_296;
         Mult_Buf[2].Weight_n = Wgt_3_296;
         Mult_Buf[3].Feature_n = FeatureBuf_297;
         Mult_Buf[3].Weight_n = Wgt_3_297;
         Mult_Buf[4].Feature_n = FeatureBuf_298;
         Mult_Buf[4].Weight_n = Wgt_3_298;
         Mult_Buf[5].Feature_n = FeatureBuf_299;
         Mult_Buf[5].Weight_n = Wgt_3_299;
         Mult_Buf[6].Feature_n = FeatureBuf_300;
         Mult_Buf[6].Weight_n = Wgt_3_300;
         Mult_Buf[7].Feature_n = FeatureBuf_301;
         Mult_Buf[7].Weight_n = Wgt_3_301;
         Mult_Buf[8].Feature_n = FeatureBuf_302;
         Mult_Buf[8].Weight_n = Wgt_3_302;
         Mult_Buf[9].Feature_n = FeatureBuf_303;
         Mult_Buf[9].Weight_n = Wgt_3_303;
         Mult_Buf[10].Feature_n = FeatureBuf_304;
         Mult_Buf[10].Weight_n = Wgt_3_304;
         Mult_Buf[11].Feature_n = FeatureBuf_305;
         Mult_Buf[11].Weight_n = Wgt_3_305;
         Mult_Buf[12].Feature_n = FeatureBuf_306;
         Mult_Buf[12].Weight_n = Wgt_3_306;
         Mult_Buf[13].Feature_n = FeatureBuf_307;
         Mult_Buf[13].Weight_n = Wgt_3_307;
         Mult_Buf[14].Feature_n = FeatureBuf_308;
         Mult_Buf[14].Weight_n = Wgt_3_308;
         Mult_Buf[15].Feature_n = FeatureBuf_309;
         Mult_Buf[15].Weight_n = Wgt_3_309;
         Mult_Buf[16].Feature_n = FeatureBuf_310;
         Mult_Buf[16].Weight_n = Wgt_3_310;
         Mult_Buf[17].Feature_n = FeatureBuf_311;
         Mult_Buf[17].Weight_n = Wgt_3_311;
         Mult_Buf[18].Feature_n = FeatureBuf_312;
         Mult_Buf[18].Weight_n = Wgt_3_312;
         Mult_Buf[19].Feature_n = FeatureBuf_313;
         Mult_Buf[19].Weight_n = Wgt_3_313;
         Mult_Buf[20].Feature_n = FeatureBuf_314;
         Mult_Buf[20].Weight_n = Wgt_3_314;
         Mult_Buf[21].Feature_n = FeatureBuf_315;
         Mult_Buf[21].Weight_n = Wgt_3_315;
         Mult_Buf[22].Feature_n = FeatureBuf_316;
         Mult_Buf[22].Weight_n = Wgt_3_316;
         Mult_Buf[23].Feature_n = FeatureBuf_317;
         Mult_Buf[23].Weight_n = Wgt_3_317;
         Mult_Buf[24].Feature_n = FeatureBuf_318;
         Mult_Buf[24].Weight_n = Wgt_3_318;
         Mult_Buf[25].Feature_n = FeatureBuf_319;
         Mult_Buf[25].Weight_n = Wgt_3_319;
         Mult_Buf[26].Feature_n = FeatureBuf_320;
         Mult_Buf[26].Weight_n = Wgt_3_320;
         Mult_Buf[27].Feature_n = FeatureBuf_321;
         Mult_Buf[27].Weight_n = Wgt_3_321;
         Mult_Buf[28].Feature_n = FeatureBuf_322;
         Mult_Buf[28].Weight_n = Wgt_3_322;
         Mult_Buf[29].Feature_n = FeatureBuf_323;
         Mult_Buf[29].Weight_n = Wgt_3_323;
         Mult_Buf[30].Feature_n = FeatureBuf_324;
         Mult_Buf[30].Weight_n = Wgt_3_324;
         Mult_Buf[31].Feature_n = FeatureBuf_325;
         Mult_Buf[31].Weight_n = Wgt_3_325;
         Mult_Buf[32].Feature_n = FeatureBuf_326;
         Mult_Buf[32].Weight_n = Wgt_3_326;
         Mult_Buf[33].Feature_n = FeatureBuf_327;
         Mult_Buf[33].Weight_n = Wgt_3_327;
         Mult_Buf[34].Feature_n = FeatureBuf_328;
         Mult_Buf[34].Weight_n = Wgt_3_328;
         Mult_Buf[35].Feature_n = FeatureBuf_329;
         Mult_Buf[35].Weight_n = Wgt_3_329;
         Mult_Buf[36].Feature_n = FeatureBuf_330;
         Mult_Buf[36].Weight_n = Wgt_3_330;
         Mult_Buf[37].Feature_n = FeatureBuf_331;
         Mult_Buf[37].Weight_n = Wgt_3_331;
         Mult_Buf[38].Feature_n = FeatureBuf_332;
         Mult_Buf[38].Weight_n = Wgt_3_332;
         Mult_Buf[39].Feature_n = FeatureBuf_333;
         Mult_Buf[39].Weight_n = Wgt_3_333;
         Mult_Buf[40].Feature_n = FeatureBuf_334;
         Mult_Buf[40].Weight_n = Wgt_3_334;
         Mult_Buf[41].Feature_n = FeatureBuf_335;
         Mult_Buf[41].Weight_n = Wgt_3_335;
         Mult_Buf[42].Feature_n = FeatureBuf_336;
         Mult_Buf[42].Weight_n = Wgt_3_336;
         Mult_Buf[43].Feature_n = FeatureBuf_337;
         Mult_Buf[43].Weight_n = Wgt_3_337;
         Mult_Buf[44].Feature_n = FeatureBuf_338;
         Mult_Buf[44].Weight_n = Wgt_3_338;
         Mult_Buf[45].Feature_n = FeatureBuf_339;
         Mult_Buf[45].Weight_n = Wgt_3_339;
         Mult_Buf[46].Feature_n = FeatureBuf_340;
         Mult_Buf[46].Weight_n = Wgt_3_340;
         Mult_Buf[47].Feature_n = FeatureBuf_341;
         Mult_Buf[47].Weight_n = Wgt_3_341;
         Mult_Buf[48].Feature_n = FeatureBuf_342;
         Mult_Buf[48].Weight_n = Wgt_3_342;
         Mult_Buf[49].Feature_n = FeatureBuf_343;
         Mult_Buf[49].Weight_n = Wgt_3_343;
         Mult_Buf[50].Feature_n = FeatureBuf_344;
         Mult_Buf[50].Weight_n = Wgt_3_344;
         Mult_Buf[51].Feature_n = FeatureBuf_345;
         Mult_Buf[51].Weight_n = Wgt_3_345;
         Mult_Buf[52].Feature_n = FeatureBuf_346;
         Mult_Buf[52].Weight_n = Wgt_3_346;
         Mult_Buf[53].Feature_n = FeatureBuf_347;
         Mult_Buf[53].Weight_n = Wgt_3_347;
         Mult_Buf[54].Feature_n = FeatureBuf_348;
         Mult_Buf[54].Weight_n = Wgt_3_348;
         Mult_Buf[55].Feature_n = FeatureBuf_349;
         Mult_Buf[55].Weight_n = Wgt_3_349;
         Mult_Buf[56].Feature_n = FeatureBuf_350;
         Mult_Buf[56].Weight_n = Wgt_3_350;
         Mult_Buf[57].Feature_n = FeatureBuf_351;
         Mult_Buf[57].Weight_n = Wgt_3_351;
         Mult_Buf[58].Feature_n = FeatureBuf_352;
         Mult_Buf[58].Weight_n = Wgt_3_352;
         Mult_Buf[59].Feature_n = FeatureBuf_353;
         Mult_Buf[59].Weight_n = Wgt_3_353;
         Mult_Buf[60].Feature_n = FeatureBuf_354;
         Mult_Buf[60].Weight_n = Wgt_3_354;
         Mult_Buf[61].Feature_n = FeatureBuf_355;
         Mult_Buf[61].Weight_n = Wgt_3_355;
         Mult_Buf[62].Feature_n = FeatureBuf_356;
         Mult_Buf[62].Weight_n = Wgt_3_356;
         Mult_Buf[63].Feature_n = FeatureBuf_357;
         Mult_Buf[63].Weight_n = Wgt_3_357;
         Mult_Buf[64].Feature_n = FeatureBuf_358;
         Mult_Buf[64].Weight_n = Wgt_3_358;
         Mult_Buf[65].Feature_n = FeatureBuf_359;
         Mult_Buf[65].Weight_n = Wgt_3_359;
         Mult_Buf[66].Feature_n = FeatureBuf_360;
         Mult_Buf[66].Weight_n = Wgt_3_360;
         Mult_Buf[67].Feature_n = FeatureBuf_361;
         Mult_Buf[67].Weight_n = Wgt_3_361;
         Mult_Buf[68].Feature_n = FeatureBuf_362;
         Mult_Buf[68].Weight_n = Wgt_3_362;
         Mult_Buf[69].Feature_n = FeatureBuf_363;
         Mult_Buf[69].Weight_n = Wgt_3_363;
         Mult_Buf[70].Feature_n = FeatureBuf_364;
         Mult_Buf[70].Weight_n = Wgt_3_364;
         Mult_Buf[71].Feature_n = FeatureBuf_365;
         Mult_Buf[71].Weight_n = Wgt_3_365;
         Mult_Buf[72].Feature_n = FeatureBuf_366;
         Mult_Buf[72].Weight_n = Wgt_3_366;
         Mult_Buf[73].Feature_n = FeatureBuf_367;
         Mult_Buf[73].Weight_n = Wgt_3_367;
         Mult_Buf[74].Feature_n = FeatureBuf_368;
         Mult_Buf[74].Weight_n = Wgt_3_368;
         Mult_Buf[75].Feature_n = FeatureBuf_369;
         Mult_Buf[75].Weight_n = Wgt_3_369;
         Mult_Buf[76].Feature_n = FeatureBuf_370;
         Mult_Buf[76].Weight_n = Wgt_3_370;
         Mult_Buf[77].Feature_n = FeatureBuf_371;
         Mult_Buf[77].Weight_n = Wgt_3_371;
         Mult_Buf[78].Feature_n = FeatureBuf_372;
         Mult_Buf[78].Weight_n = Wgt_3_372;
         Mult_Buf[79].Feature_n = FeatureBuf_373;
         Mult_Buf[79].Weight_n = Wgt_3_373;
         Mult_Buf[80].Feature_n = FeatureBuf_374;
         Mult_Buf[80].Weight_n = Wgt_3_374;
         Mult_Buf[81].Feature_n = FeatureBuf_375;
         Mult_Buf[81].Weight_n = Wgt_3_375;
         Mult_Buf[82].Feature_n = FeatureBuf_376;
         Mult_Buf[82].Weight_n = Wgt_3_376;
         Mult_Buf[83].Feature_n = FeatureBuf_377;
         Mult_Buf[83].Weight_n = Wgt_3_377;
         Mult_Buf[84].Feature_n = FeatureBuf_378;
         Mult_Buf[84].Weight_n = Wgt_3_378;
         Mult_Buf[85].Feature_n = FeatureBuf_379;
         Mult_Buf[85].Weight_n = Wgt_3_379;
         Mult_Buf[86].Feature_n = FeatureBuf_380;
         Mult_Buf[86].Weight_n = Wgt_3_380;
         Mult_Buf[87].Feature_n = FeatureBuf_381;
         Mult_Buf[87].Weight_n = Wgt_3_381;
         Mult_Buf[88].Feature_n = FeatureBuf_382;
         Mult_Buf[88].Weight_n = Wgt_3_382;
         Mult_Buf[89].Feature_n = FeatureBuf_383;
         Mult_Buf[89].Weight_n = Wgt_3_383;
         Mult_Buf[90].Feature_n = FeatureBuf_384;
         Mult_Buf[90].Weight_n = Wgt_3_384;
         Mult_Buf[91].Feature_n = FeatureBuf_385;
         Mult_Buf[91].Weight_n = Wgt_3_385;
         Mult_Buf[92].Feature_n = FeatureBuf_386;
         Mult_Buf[92].Weight_n = Wgt_3_386;
         Mult_Buf[93].Feature_n = FeatureBuf_387;
         Mult_Buf[93].Weight_n = Wgt_3_387;
         Mult_Buf[94].Feature_n = FeatureBuf_388;
         Mult_Buf[94].Weight_n = Wgt_3_388;
         Mult_Buf[95].Feature_n = FeatureBuf_389;
         Mult_Buf[95].Weight_n = Wgt_3_389;
         Mult_Buf[96].Feature_n = FeatureBuf_390;
         Mult_Buf[96].Weight_n = Wgt_3_390;
         Mult_Buf[97].Feature_n = FeatureBuf_391;
         Mult_Buf[97].Weight_n = Wgt_3_391;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     //Collect Partial result form Adder
         Res_0_5_n = Part_Res;
     end
    30:begin
     nxt_state = 31;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_392;
         Mult_Buf[0].Weight_n = Wgt_3_392;
         Mult_Buf[1].Feature_n = FeatureBuf_393;
         Mult_Buf[1].Weight_n = Wgt_3_393;
         Mult_Buf[2].Feature_n = FeatureBuf_394;
         Mult_Buf[2].Weight_n = Wgt_3_394;
         Mult_Buf[3].Feature_n = FeatureBuf_395;
         Mult_Buf[3].Weight_n = Wgt_3_395;
         Mult_Buf[4].Feature_n = FeatureBuf_396;
         Mult_Buf[4].Weight_n = Wgt_3_396;
         Mult_Buf[5].Feature_n = FeatureBuf_397;
         Mult_Buf[5].Weight_n = Wgt_3_397;
         Mult_Buf[6].Feature_n = FeatureBuf_398;
         Mult_Buf[6].Weight_n = Wgt_3_398;
         Mult_Buf[7].Feature_n = FeatureBuf_399;
         Mult_Buf[7].Weight_n = Wgt_3_399;
         Mult_Buf[8].Feature_n = FeatureBuf_400;
         Mult_Buf[8].Weight_n = Wgt_3_400;
         Mult_Buf[9].Feature_n = FeatureBuf_401;
         Mult_Buf[9].Weight_n = Wgt_3_401;
         Mult_Buf[10].Feature_n = FeatureBuf_402;
         Mult_Buf[10].Weight_n = Wgt_3_402;
         Mult_Buf[11].Feature_n = FeatureBuf_403;
         Mult_Buf[11].Weight_n = Wgt_3_403;
         Mult_Buf[12].Feature_n = FeatureBuf_404;
         Mult_Buf[12].Weight_n = Wgt_3_404;
         Mult_Buf[13].Feature_n = FeatureBuf_405;
         Mult_Buf[13].Weight_n = Wgt_3_405;
         Mult_Buf[14].Feature_n = FeatureBuf_406;
         Mult_Buf[14].Weight_n = Wgt_3_406;
         Mult_Buf[15].Feature_n = FeatureBuf_407;
         Mult_Buf[15].Weight_n = Wgt_3_407;
         Mult_Buf[16].Feature_n = FeatureBuf_408;
         Mult_Buf[16].Weight_n = Wgt_3_408;
         Mult_Buf[17].Feature_n = FeatureBuf_409;
         Mult_Buf[17].Weight_n = Wgt_3_409;
         Mult_Buf[18].Feature_n = FeatureBuf_410;
         Mult_Buf[18].Weight_n = Wgt_3_410;
         Mult_Buf[19].Feature_n = FeatureBuf_411;
         Mult_Buf[19].Weight_n = Wgt_3_411;
         Mult_Buf[20].Feature_n = FeatureBuf_412;
         Mult_Buf[20].Weight_n = Wgt_3_412;
         Mult_Buf[21].Feature_n = FeatureBuf_413;
         Mult_Buf[21].Weight_n = Wgt_3_413;
         Mult_Buf[22].Feature_n = FeatureBuf_414;
         Mult_Buf[22].Weight_n = Wgt_3_414;
         Mult_Buf[23].Feature_n = FeatureBuf_415;
         Mult_Buf[23].Weight_n = Wgt_3_415;
         Mult_Buf[24].Feature_n = FeatureBuf_416;
         Mult_Buf[24].Weight_n = Wgt_3_416;
         Mult_Buf[25].Feature_n = FeatureBuf_417;
         Mult_Buf[25].Weight_n = Wgt_3_417;
         Mult_Buf[26].Feature_n = FeatureBuf_418;
         Mult_Buf[26].Weight_n = Wgt_3_418;
         Mult_Buf[27].Feature_n = FeatureBuf_419;
         Mult_Buf[27].Weight_n = Wgt_3_419;
         Mult_Buf[28].Feature_n = FeatureBuf_420;
         Mult_Buf[28].Weight_n = Wgt_3_420;
         Mult_Buf[29].Feature_n = FeatureBuf_421;
         Mult_Buf[29].Weight_n = Wgt_3_421;
         Mult_Buf[30].Feature_n = FeatureBuf_422;
         Mult_Buf[30].Weight_n = Wgt_3_422;
         Mult_Buf[31].Feature_n = FeatureBuf_423;
         Mult_Buf[31].Weight_n = Wgt_3_423;
         Mult_Buf[32].Feature_n = FeatureBuf_424;
         Mult_Buf[32].Weight_n = Wgt_3_424;
         Mult_Buf[33].Feature_n = FeatureBuf_425;
         Mult_Buf[33].Weight_n = Wgt_3_425;
         Mult_Buf[34].Feature_n = FeatureBuf_426;
         Mult_Buf[34].Weight_n = Wgt_3_426;
         Mult_Buf[35].Feature_n = FeatureBuf_427;
         Mult_Buf[35].Weight_n = Wgt_3_427;
         Mult_Buf[36].Feature_n = FeatureBuf_428;
         Mult_Buf[36].Weight_n = Wgt_3_428;
         Mult_Buf[37].Feature_n = FeatureBuf_429;
         Mult_Buf[37].Weight_n = Wgt_3_429;
         Mult_Buf[38].Feature_n = FeatureBuf_430;
         Mult_Buf[38].Weight_n = Wgt_3_430;
         Mult_Buf[39].Feature_n = FeatureBuf_431;
         Mult_Buf[39].Weight_n = Wgt_3_431;
         Mult_Buf[40].Feature_n = FeatureBuf_432;
         Mult_Buf[40].Weight_n = Wgt_3_432;
         Mult_Buf[41].Feature_n = FeatureBuf_433;
         Mult_Buf[41].Weight_n = Wgt_3_433;
         Mult_Buf[42].Feature_n = FeatureBuf_434;
         Mult_Buf[42].Weight_n = Wgt_3_434;
         Mult_Buf[43].Feature_n = FeatureBuf_435;
         Mult_Buf[43].Weight_n = Wgt_3_435;
         Mult_Buf[44].Feature_n = FeatureBuf_436;
         Mult_Buf[44].Weight_n = Wgt_3_436;
         Mult_Buf[45].Feature_n = FeatureBuf_437;
         Mult_Buf[45].Weight_n = Wgt_3_437;
         Mult_Buf[46].Feature_n = FeatureBuf_438;
         Mult_Buf[46].Weight_n = Wgt_3_438;
         Mult_Buf[47].Feature_n = FeatureBuf_439;
         Mult_Buf[47].Weight_n = Wgt_3_439;
         Mult_Buf[48].Feature_n = FeatureBuf_440;
         Mult_Buf[48].Weight_n = Wgt_3_440;
         Mult_Buf[49].Feature_n = FeatureBuf_441;
         Mult_Buf[49].Weight_n = Wgt_3_441;
         Mult_Buf[50].Feature_n = FeatureBuf_442;
         Mult_Buf[50].Weight_n = Wgt_3_442;
         Mult_Buf[51].Feature_n = FeatureBuf_443;
         Mult_Buf[51].Weight_n = Wgt_3_443;
         Mult_Buf[52].Feature_n = FeatureBuf_444;
         Mult_Buf[52].Weight_n = Wgt_3_444;
         Mult_Buf[53].Feature_n = FeatureBuf_445;
         Mult_Buf[53].Weight_n = Wgt_3_445;
         Mult_Buf[54].Feature_n = FeatureBuf_446;
         Mult_Buf[54].Weight_n = Wgt_3_446;
         Mult_Buf[55].Feature_n = FeatureBuf_447;
         Mult_Buf[55].Weight_n = Wgt_3_447;
         Mult_Buf[56].Feature_n = FeatureBuf_448;
         Mult_Buf[56].Weight_n = Wgt_3_448;
         Mult_Buf[57].Feature_n = FeatureBuf_449;
         Mult_Buf[57].Weight_n = Wgt_3_449;
         Mult_Buf[58].Feature_n = FeatureBuf_450;
         Mult_Buf[58].Weight_n = Wgt_3_450;
         Mult_Buf[59].Feature_n = FeatureBuf_451;
         Mult_Buf[59].Weight_n = Wgt_3_451;
         Mult_Buf[60].Feature_n = FeatureBuf_452;
         Mult_Buf[60].Weight_n = Wgt_3_452;
         Mult_Buf[61].Feature_n = FeatureBuf_453;
         Mult_Buf[61].Weight_n = Wgt_3_453;
         Mult_Buf[62].Feature_n = FeatureBuf_454;
         Mult_Buf[62].Weight_n = Wgt_3_454;
         Mult_Buf[63].Feature_n = FeatureBuf_455;
         Mult_Buf[63].Weight_n = Wgt_3_455;
         Mult_Buf[64].Feature_n = FeatureBuf_456;
         Mult_Buf[64].Weight_n = Wgt_3_456;
         Mult_Buf[65].Feature_n = FeatureBuf_457;
         Mult_Buf[65].Weight_n = Wgt_3_457;
         Mult_Buf[66].Feature_n = FeatureBuf_458;
         Mult_Buf[66].Weight_n = Wgt_3_458;
         Mult_Buf[67].Feature_n = FeatureBuf_459;
         Mult_Buf[67].Weight_n = Wgt_3_459;
         Mult_Buf[68].Feature_n = FeatureBuf_460;
         Mult_Buf[68].Weight_n = Wgt_3_460;
         Mult_Buf[69].Feature_n = FeatureBuf_461;
         Mult_Buf[69].Weight_n = Wgt_3_461;
         Mult_Buf[70].Feature_n = FeatureBuf_462;
         Mult_Buf[70].Weight_n = Wgt_3_462;
         Mult_Buf[71].Feature_n = FeatureBuf_463;
         Mult_Buf[71].Weight_n = Wgt_3_463;
         Mult_Buf[72].Feature_n = FeatureBuf_464;
         Mult_Buf[72].Weight_n = Wgt_3_464;
         Mult_Buf[73].Feature_n = FeatureBuf_465;
         Mult_Buf[73].Weight_n = Wgt_3_465;
         Mult_Buf[74].Feature_n = FeatureBuf_466;
         Mult_Buf[74].Weight_n = Wgt_3_466;
         Mult_Buf[75].Feature_n = FeatureBuf_467;
         Mult_Buf[75].Weight_n = Wgt_3_467;
         Mult_Buf[76].Feature_n = FeatureBuf_468;
         Mult_Buf[76].Weight_n = Wgt_3_468;
         Mult_Buf[77].Feature_n = FeatureBuf_469;
         Mult_Buf[77].Weight_n = Wgt_3_469;
         Mult_Buf[78].Feature_n = FeatureBuf_470;
         Mult_Buf[78].Weight_n = Wgt_3_470;
         Mult_Buf[79].Feature_n = FeatureBuf_471;
         Mult_Buf[79].Weight_n = Wgt_3_471;
         Mult_Buf[80].Feature_n = FeatureBuf_472;
         Mult_Buf[80].Weight_n = Wgt_3_472;
         Mult_Buf[81].Feature_n = FeatureBuf_473;
         Mult_Buf[81].Weight_n = Wgt_3_473;
         Mult_Buf[82].Feature_n = FeatureBuf_474;
         Mult_Buf[82].Weight_n = Wgt_3_474;
         Mult_Buf[83].Feature_n = FeatureBuf_475;
         Mult_Buf[83].Weight_n = Wgt_3_475;
         Mult_Buf[84].Feature_n = FeatureBuf_476;
         Mult_Buf[84].Weight_n = Wgt_3_476;
         Mult_Buf[85].Feature_n = FeatureBuf_477;
         Mult_Buf[85].Weight_n = Wgt_3_477;
         Mult_Buf[86].Feature_n = FeatureBuf_478;
         Mult_Buf[86].Weight_n = Wgt_3_478;
         Mult_Buf[87].Feature_n = FeatureBuf_479;
         Mult_Buf[87].Weight_n = Wgt_3_479;
         Mult_Buf[88].Feature_n = FeatureBuf_480;
         Mult_Buf[88].Weight_n = Wgt_3_480;
         Mult_Buf[89].Feature_n = FeatureBuf_481;
         Mult_Buf[89].Weight_n = Wgt_3_481;
         Mult_Buf[90].Feature_n = FeatureBuf_482;
         Mult_Buf[90].Weight_n = Wgt_3_482;
         Mult_Buf[91].Feature_n = FeatureBuf_483;
         Mult_Buf[91].Weight_n = Wgt_3_483;
         Mult_Buf[92].Feature_n = FeatureBuf_484;
         Mult_Buf[92].Weight_n = Wgt_3_484;
         Mult_Buf[93].Feature_n = FeatureBuf_485;
         Mult_Buf[93].Weight_n = Wgt_3_485;
         Mult_Buf[94].Feature_n = FeatureBuf_486;
         Mult_Buf[94].Weight_n = Wgt_3_486;
         Mult_Buf[95].Feature_n = FeatureBuf_487;
         Mult_Buf[95].Weight_n = Wgt_3_487;
         Mult_Buf[96].Feature_n = FeatureBuf_488;
         Mult_Buf[96].Weight_n = Wgt_3_488;
         Mult_Buf[97].Feature_n = FeatureBuf_489;
         Mult_Buf[97].Weight_n = Wgt_3_489;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     //Collect Partial result form Adder
         Res_0_6_n = Part_Res;
     end
    31:begin
     nxt_state = 32;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_490;
         Mult_Buf[0].Weight_n = Wgt_3_490;
         Mult_Buf[1].Feature_n = FeatureBuf_491;
         Mult_Buf[1].Weight_n = Wgt_3_491;
         Mult_Buf[2].Feature_n = FeatureBuf_492;
         Mult_Buf[2].Weight_n = Wgt_3_492;
         Mult_Buf[3].Feature_n = FeatureBuf_493;
         Mult_Buf[3].Weight_n = Wgt_3_493;
         Mult_Buf[4].Feature_n = FeatureBuf_494;
         Mult_Buf[4].Weight_n = Wgt_3_494;
         Mult_Buf[5].Feature_n = FeatureBuf_495;
         Mult_Buf[5].Weight_n = Wgt_3_495;
         Mult_Buf[6].Feature_n = FeatureBuf_496;
         Mult_Buf[6].Weight_n = Wgt_3_496;
         Mult_Buf[7].Feature_n = FeatureBuf_497;
         Mult_Buf[7].Weight_n = Wgt_3_497;
         Mult_Buf[8].Feature_n = FeatureBuf_498;
         Mult_Buf[8].Weight_n = Wgt_3_498;
         Mult_Buf[9].Feature_n = FeatureBuf_499;
         Mult_Buf[9].Weight_n = Wgt_3_499;
         Mult_Buf[10].Feature_n = FeatureBuf_500;
         Mult_Buf[10].Weight_n = Wgt_3_500;
         Mult_Buf[11].Feature_n = FeatureBuf_501;
         Mult_Buf[11].Weight_n = Wgt_3_501;
         Mult_Buf[12].Feature_n = FeatureBuf_502;
         Mult_Buf[12].Weight_n = Wgt_3_502;
         Mult_Buf[13].Feature_n = FeatureBuf_503;
         Mult_Buf[13].Weight_n = Wgt_3_503;
         Mult_Buf[14].Feature_n = FeatureBuf_504;
         Mult_Buf[14].Weight_n = Wgt_3_504;
         Mult_Buf[15].Feature_n = FeatureBuf_505;
         Mult_Buf[15].Weight_n = Wgt_3_505;
         Mult_Buf[16].Feature_n = FeatureBuf_506;
         Mult_Buf[16].Weight_n = Wgt_3_506;
         Mult_Buf[17].Feature_n = FeatureBuf_507;
         Mult_Buf[17].Weight_n = Wgt_3_507;
         Mult_Buf[18].Feature_n = FeatureBuf_508;
         Mult_Buf[18].Weight_n = Wgt_3_508;
         Mult_Buf[19].Feature_n = FeatureBuf_509;
         Mult_Buf[19].Weight_n = Wgt_3_509;
         Mult_Buf[20].Feature_n = FeatureBuf_510;
         Mult_Buf[20].Weight_n = Wgt_3_510;
         Mult_Buf[21].Feature_n = FeatureBuf_511;
         Mult_Buf[21].Weight_n = Wgt_3_511;
         Mult_Buf[22].Feature_n = FeatureBuf_512;
         Mult_Buf[22].Weight_n = Wgt_3_512;
         Mult_Buf[23].Feature_n = FeatureBuf_513;
         Mult_Buf[23].Weight_n = Wgt_3_513;
         Mult_Buf[24].Feature_n = FeatureBuf_514;
         Mult_Buf[24].Weight_n = Wgt_3_514;
         Mult_Buf[25].Feature_n = FeatureBuf_515;
         Mult_Buf[25].Weight_n = Wgt_3_515;
         Mult_Buf[26].Feature_n = FeatureBuf_516;
         Mult_Buf[26].Weight_n = Wgt_3_516;
         Mult_Buf[27].Feature_n = FeatureBuf_517;
         Mult_Buf[27].Weight_n = Wgt_3_517;
         Mult_Buf[28].Feature_n = FeatureBuf_518;
         Mult_Buf[28].Weight_n = Wgt_3_518;
         Mult_Buf[29].Feature_n = FeatureBuf_519;
         Mult_Buf[29].Weight_n = Wgt_3_519;
         Mult_Buf[30].Feature_n = FeatureBuf_520;
         Mult_Buf[30].Weight_n = Wgt_3_520;
         Mult_Buf[31].Feature_n = FeatureBuf_521;
         Mult_Buf[31].Weight_n = Wgt_3_521;
         Mult_Buf[32].Feature_n = FeatureBuf_522;
         Mult_Buf[32].Weight_n = Wgt_3_522;
         Mult_Buf[33].Feature_n = FeatureBuf_523;
         Mult_Buf[33].Weight_n = Wgt_3_523;
         Mult_Buf[34].Feature_n = FeatureBuf_524;
         Mult_Buf[34].Weight_n = Wgt_3_524;
         Mult_Buf[35].Feature_n = FeatureBuf_525;
         Mult_Buf[35].Weight_n = Wgt_3_525;
         Mult_Buf[36].Feature_n = FeatureBuf_526;
         Mult_Buf[36].Weight_n = Wgt_3_526;
         Mult_Buf[37].Feature_n = FeatureBuf_527;
         Mult_Buf[37].Weight_n = Wgt_3_527;
         Mult_Buf[38].Feature_n = FeatureBuf_528;
         Mult_Buf[38].Weight_n = Wgt_3_528;
         Mult_Buf[39].Feature_n = FeatureBuf_529;
         Mult_Buf[39].Weight_n = Wgt_3_529;
         Mult_Buf[40].Feature_n = FeatureBuf_530;
         Mult_Buf[40].Weight_n = Wgt_3_530;
         Mult_Buf[41].Feature_n = FeatureBuf_531;
         Mult_Buf[41].Weight_n = Wgt_3_531;
         Mult_Buf[42].Feature_n = FeatureBuf_532;
         Mult_Buf[42].Weight_n = Wgt_3_532;
         Mult_Buf[43].Feature_n = FeatureBuf_533;
         Mult_Buf[43].Weight_n = Wgt_3_533;
         Mult_Buf[44].Feature_n = FeatureBuf_534;
         Mult_Buf[44].Weight_n = Wgt_3_534;
         Mult_Buf[45].Feature_n = FeatureBuf_535;
         Mult_Buf[45].Weight_n = Wgt_3_535;
         Mult_Buf[46].Feature_n = FeatureBuf_536;
         Mult_Buf[46].Weight_n = Wgt_3_536;
         Mult_Buf[47].Feature_n = FeatureBuf_537;
         Mult_Buf[47].Weight_n = Wgt_3_537;
         Mult_Buf[48].Feature_n = FeatureBuf_538;
         Mult_Buf[48].Weight_n = Wgt_3_538;
         Mult_Buf[49].Feature_n = FeatureBuf_539;
         Mult_Buf[49].Weight_n = Wgt_3_539;
         Mult_Buf[50].Feature_n = FeatureBuf_540;
         Mult_Buf[50].Weight_n = Wgt_3_540;
         Mult_Buf[51].Feature_n = FeatureBuf_541;
         Mult_Buf[51].Weight_n = Wgt_3_541;
         Mult_Buf[52].Feature_n = FeatureBuf_542;
         Mult_Buf[52].Weight_n = Wgt_3_542;
         Mult_Buf[53].Feature_n = FeatureBuf_543;
         Mult_Buf[53].Weight_n = Wgt_3_543;
         Mult_Buf[54].Feature_n = FeatureBuf_544;
         Mult_Buf[54].Weight_n = Wgt_3_544;
         Mult_Buf[55].Feature_n = FeatureBuf_545;
         Mult_Buf[55].Weight_n = Wgt_3_545;
         Mult_Buf[56].Feature_n = FeatureBuf_546;
         Mult_Buf[56].Weight_n = Wgt_3_546;
         Mult_Buf[57].Feature_n = FeatureBuf_547;
         Mult_Buf[57].Weight_n = Wgt_3_547;
         Mult_Buf[58].Feature_n = FeatureBuf_548;
         Mult_Buf[58].Weight_n = Wgt_3_548;
         Mult_Buf[59].Feature_n = FeatureBuf_549;
         Mult_Buf[59].Weight_n = Wgt_3_549;
         Mult_Buf[60].Feature_n = FeatureBuf_550;
         Mult_Buf[60].Weight_n = Wgt_3_550;
         Mult_Buf[61].Feature_n = FeatureBuf_551;
         Mult_Buf[61].Weight_n = Wgt_3_551;
         Mult_Buf[62].Feature_n = FeatureBuf_552;
         Mult_Buf[62].Weight_n = Wgt_3_552;
         Mult_Buf[63].Feature_n = FeatureBuf_553;
         Mult_Buf[63].Weight_n = Wgt_3_553;
         Mult_Buf[64].Feature_n = FeatureBuf_554;
         Mult_Buf[64].Weight_n = Wgt_3_554;
         Mult_Buf[65].Feature_n = FeatureBuf_555;
         Mult_Buf[65].Weight_n = Wgt_3_555;
         Mult_Buf[66].Feature_n = FeatureBuf_556;
         Mult_Buf[66].Weight_n = Wgt_3_556;
         Mult_Buf[67].Feature_n = FeatureBuf_557;
         Mult_Buf[67].Weight_n = Wgt_3_557;
         Mult_Buf[68].Feature_n = FeatureBuf_558;
         Mult_Buf[68].Weight_n = Wgt_3_558;
         Mult_Buf[69].Feature_n = FeatureBuf_559;
         Mult_Buf[69].Weight_n = Wgt_3_559;
         Mult_Buf[70].Feature_n = FeatureBuf_560;
         Mult_Buf[70].Weight_n = Wgt_3_560;
         Mult_Buf[71].Feature_n = FeatureBuf_561;
         Mult_Buf[71].Weight_n = Wgt_3_561;
         Mult_Buf[72].Feature_n = FeatureBuf_562;
         Mult_Buf[72].Weight_n = Wgt_3_562;
         Mult_Buf[73].Feature_n = FeatureBuf_563;
         Mult_Buf[73].Weight_n = Wgt_3_563;
         Mult_Buf[74].Feature_n = FeatureBuf_564;
         Mult_Buf[74].Weight_n = Wgt_3_564;
         Mult_Buf[75].Feature_n = FeatureBuf_565;
         Mult_Buf[75].Weight_n = Wgt_3_565;
         Mult_Buf[76].Feature_n = FeatureBuf_566;
         Mult_Buf[76].Weight_n = Wgt_3_566;
         Mult_Buf[77].Feature_n = FeatureBuf_567;
         Mult_Buf[77].Weight_n = Wgt_3_567;
         Mult_Buf[78].Feature_n = FeatureBuf_568;
         Mult_Buf[78].Weight_n = Wgt_3_568;
         Mult_Buf[79].Feature_n = FeatureBuf_569;
         Mult_Buf[79].Weight_n = Wgt_3_569;
         Mult_Buf[80].Feature_n = FeatureBuf_570;
         Mult_Buf[80].Weight_n = Wgt_3_570;
         Mult_Buf[81].Feature_n = FeatureBuf_571;
         Mult_Buf[81].Weight_n = Wgt_3_571;
         Mult_Buf[82].Feature_n = FeatureBuf_572;
         Mult_Buf[82].Weight_n = Wgt_3_572;
         Mult_Buf[83].Feature_n = FeatureBuf_573;
         Mult_Buf[83].Weight_n = Wgt_3_573;
         Mult_Buf[84].Feature_n = FeatureBuf_574;
         Mult_Buf[84].Weight_n = Wgt_3_574;
         Mult_Buf[85].Feature_n = FeatureBuf_575;
         Mult_Buf[85].Weight_n = Wgt_3_575;
         Mult_Buf[86].Feature_n = FeatureBuf_576;
         Mult_Buf[86].Weight_n = Wgt_3_576;
         Mult_Buf[87].Feature_n = FeatureBuf_577;
         Mult_Buf[87].Weight_n = Wgt_3_577;
         Mult_Buf[88].Feature_n = FeatureBuf_578;
         Mult_Buf[88].Weight_n = Wgt_3_578;
         Mult_Buf[89].Feature_n = FeatureBuf_579;
         Mult_Buf[89].Weight_n = Wgt_3_579;
         Mult_Buf[90].Feature_n = FeatureBuf_580;
         Mult_Buf[90].Weight_n = Wgt_3_580;
         Mult_Buf[91].Feature_n = FeatureBuf_581;
         Mult_Buf[91].Weight_n = Wgt_3_581;
         Mult_Buf[92].Feature_n = FeatureBuf_582;
         Mult_Buf[92].Weight_n = Wgt_3_582;
         Mult_Buf[93].Feature_n = FeatureBuf_583;
         Mult_Buf[93].Weight_n = Wgt_3_583;
         Mult_Buf[94].Feature_n = FeatureBuf_584;
         Mult_Buf[94].Weight_n = Wgt_3_584;
         Mult_Buf[95].Feature_n = FeatureBuf_585;
         Mult_Buf[95].Weight_n = Wgt_3_585;
         Mult_Buf[96].Feature_n = FeatureBuf_586;
         Mult_Buf[96].Weight_n = Wgt_3_586;
         Mult_Buf[97].Feature_n = FeatureBuf_587;
         Mult_Buf[97].Weight_n = Wgt_3_587;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     //Collect Partial result form Adder
         Res_0_7_n = Part_Res;
     //Feed to final Adder
         A1 = Part_Res;
         A2 = Res_0_6_n;
         A3 = Res_0_5_n;
         A4 = Res_0_4_n;
         A5 = Res_0_3_n;
         A6 = Res_0_2_n;
         A7 = Res_0_1_n;
         A8 = Res_0_0_n;
     end
    32:begin
     nxt_state = 33;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_588;
         Mult_Buf[0].Weight_n = Wgt_3_588;
         Mult_Buf[1].Feature_n = FeatureBuf_589;
         Mult_Buf[1].Weight_n = Wgt_3_589;
         Mult_Buf[2].Feature_n = FeatureBuf_590;
         Mult_Buf[2].Weight_n = Wgt_3_590;
         Mult_Buf[3].Feature_n = FeatureBuf_591;
         Mult_Buf[3].Weight_n = Wgt_3_591;
         Mult_Buf[4].Feature_n = FeatureBuf_592;
         Mult_Buf[4].Weight_n = Wgt_3_592;
         Mult_Buf[5].Feature_n = FeatureBuf_593;
         Mult_Buf[5].Weight_n = Wgt_3_593;
         Mult_Buf[6].Feature_n = FeatureBuf_594;
         Mult_Buf[6].Weight_n = Wgt_3_594;
         Mult_Buf[7].Feature_n = FeatureBuf_595;
         Mult_Buf[7].Weight_n = Wgt_3_595;
         Mult_Buf[8].Feature_n = FeatureBuf_596;
         Mult_Buf[8].Weight_n = Wgt_3_596;
         Mult_Buf[9].Feature_n = FeatureBuf_597;
         Mult_Buf[9].Weight_n = Wgt_3_597;
         Mult_Buf[10].Feature_n = FeatureBuf_598;
         Mult_Buf[10].Weight_n = Wgt_3_598;
         Mult_Buf[11].Feature_n = FeatureBuf_599;
         Mult_Buf[11].Weight_n = Wgt_3_599;
         Mult_Buf[12].Feature_n = FeatureBuf_600;
         Mult_Buf[12].Weight_n = Wgt_3_600;
         Mult_Buf[13].Feature_n = FeatureBuf_601;
         Mult_Buf[13].Weight_n = Wgt_3_601;
         Mult_Buf[14].Feature_n = FeatureBuf_602;
         Mult_Buf[14].Weight_n = Wgt_3_602;
         Mult_Buf[15].Feature_n = FeatureBuf_603;
         Mult_Buf[15].Weight_n = Wgt_3_603;
         Mult_Buf[16].Feature_n = FeatureBuf_604;
         Mult_Buf[16].Weight_n = Wgt_3_604;
         Mult_Buf[17].Feature_n = FeatureBuf_605;
         Mult_Buf[17].Weight_n = Wgt_3_605;
         Mult_Buf[18].Feature_n = FeatureBuf_606;
         Mult_Buf[18].Weight_n = Wgt_3_606;
         Mult_Buf[19].Feature_n = FeatureBuf_607;
         Mult_Buf[19].Weight_n = Wgt_3_607;
         Mult_Buf[20].Feature_n = FeatureBuf_608;
         Mult_Buf[20].Weight_n = Wgt_3_608;
         Mult_Buf[21].Feature_n = FeatureBuf_609;
         Mult_Buf[21].Weight_n = Wgt_3_609;
         Mult_Buf[22].Feature_n = FeatureBuf_610;
         Mult_Buf[22].Weight_n = Wgt_3_610;
         Mult_Buf[23].Feature_n = FeatureBuf_611;
         Mult_Buf[23].Weight_n = Wgt_3_611;
         Mult_Buf[24].Feature_n = FeatureBuf_612;
         Mult_Buf[24].Weight_n = Wgt_3_612;
         Mult_Buf[25].Feature_n = FeatureBuf_613;
         Mult_Buf[25].Weight_n = Wgt_3_613;
         Mult_Buf[26].Feature_n = FeatureBuf_614;
         Mult_Buf[26].Weight_n = Wgt_3_614;
         Mult_Buf[27].Feature_n = FeatureBuf_615;
         Mult_Buf[27].Weight_n = Wgt_3_615;
         Mult_Buf[28].Feature_n = FeatureBuf_616;
         Mult_Buf[28].Weight_n = Wgt_3_616;
         Mult_Buf[29].Feature_n = FeatureBuf_617;
         Mult_Buf[29].Weight_n = Wgt_3_617;
         Mult_Buf[30].Feature_n = FeatureBuf_618;
         Mult_Buf[30].Weight_n = Wgt_3_618;
         Mult_Buf[31].Feature_n = FeatureBuf_619;
         Mult_Buf[31].Weight_n = Wgt_3_619;
         Mult_Buf[32].Feature_n = FeatureBuf_620;
         Mult_Buf[32].Weight_n = Wgt_3_620;
         Mult_Buf[33].Feature_n = FeatureBuf_621;
         Mult_Buf[33].Weight_n = Wgt_3_621;
         Mult_Buf[34].Feature_n = FeatureBuf_622;
         Mult_Buf[34].Weight_n = Wgt_3_622;
         Mult_Buf[35].Feature_n = FeatureBuf_623;
         Mult_Buf[35].Weight_n = Wgt_3_623;
         Mult_Buf[36].Feature_n = FeatureBuf_624;
         Mult_Buf[36].Weight_n = Wgt_3_624;
         Mult_Buf[37].Feature_n = FeatureBuf_625;
         Mult_Buf[37].Weight_n = Wgt_3_625;
         Mult_Buf[38].Feature_n = FeatureBuf_626;
         Mult_Buf[38].Weight_n = Wgt_3_626;
         Mult_Buf[39].Feature_n = FeatureBuf_627;
         Mult_Buf[39].Weight_n = Wgt_3_627;
         Mult_Buf[40].Feature_n = FeatureBuf_628;
         Mult_Buf[40].Weight_n = Wgt_3_628;
         Mult_Buf[41].Feature_n = FeatureBuf_629;
         Mult_Buf[41].Weight_n = Wgt_3_629;
         Mult_Buf[42].Feature_n = FeatureBuf_630;
         Mult_Buf[42].Weight_n = Wgt_3_630;
         Mult_Buf[43].Feature_n = FeatureBuf_631;
         Mult_Buf[43].Weight_n = Wgt_3_631;
         Mult_Buf[44].Feature_n = FeatureBuf_632;
         Mult_Buf[44].Weight_n = Wgt_3_632;
         Mult_Buf[45].Feature_n = FeatureBuf_633;
         Mult_Buf[45].Weight_n = Wgt_3_633;
         Mult_Buf[46].Feature_n = FeatureBuf_634;
         Mult_Buf[46].Weight_n = Wgt_3_634;
         Mult_Buf[47].Feature_n = FeatureBuf_635;
         Mult_Buf[47].Weight_n = Wgt_3_635;
         Mult_Buf[48].Feature_n = FeatureBuf_636;
         Mult_Buf[48].Weight_n = Wgt_3_636;
         Mult_Buf[49].Feature_n = FeatureBuf_637;
         Mult_Buf[49].Weight_n = Wgt_3_637;
         Mult_Buf[50].Feature_n = FeatureBuf_638;
         Mult_Buf[50].Weight_n = Wgt_3_638;
         Mult_Buf[51].Feature_n = FeatureBuf_639;
         Mult_Buf[51].Weight_n = Wgt_3_639;
         Mult_Buf[52].Feature_n = FeatureBuf_640;
         Mult_Buf[52].Weight_n = Wgt_3_640;
         Mult_Buf[53].Feature_n = FeatureBuf_641;
         Mult_Buf[53].Weight_n = Wgt_3_641;
         Mult_Buf[54].Feature_n = FeatureBuf_642;
         Mult_Buf[54].Weight_n = Wgt_3_642;
         Mult_Buf[55].Feature_n = FeatureBuf_643;
         Mult_Buf[55].Weight_n = Wgt_3_643;
         Mult_Buf[56].Feature_n = FeatureBuf_644;
         Mult_Buf[56].Weight_n = Wgt_3_644;
         Mult_Buf[57].Feature_n = FeatureBuf_645;
         Mult_Buf[57].Weight_n = Wgt_3_645;
         Mult_Buf[58].Feature_n = FeatureBuf_646;
         Mult_Buf[58].Weight_n = Wgt_3_646;
         Mult_Buf[59].Feature_n = FeatureBuf_647;
         Mult_Buf[59].Weight_n = Wgt_3_647;
         Mult_Buf[60].Feature_n = FeatureBuf_648;
         Mult_Buf[60].Weight_n = Wgt_3_648;
         Mult_Buf[61].Feature_n = FeatureBuf_649;
         Mult_Buf[61].Weight_n = Wgt_3_649;
         Mult_Buf[62].Feature_n = FeatureBuf_650;
         Mult_Buf[62].Weight_n = Wgt_3_650;
         Mult_Buf[63].Feature_n = FeatureBuf_651;
         Mult_Buf[63].Weight_n = Wgt_3_651;
         Mult_Buf[64].Feature_n = FeatureBuf_652;
         Mult_Buf[64].Weight_n = Wgt_3_652;
         Mult_Buf[65].Feature_n = FeatureBuf_653;
         Mult_Buf[65].Weight_n = Wgt_3_653;
         Mult_Buf[66].Feature_n = FeatureBuf_654;
         Mult_Buf[66].Weight_n = Wgt_3_654;
         Mult_Buf[67].Feature_n = FeatureBuf_655;
         Mult_Buf[67].Weight_n = Wgt_3_655;
         Mult_Buf[68].Feature_n = FeatureBuf_656;
         Mult_Buf[68].Weight_n = Wgt_3_656;
         Mult_Buf[69].Feature_n = FeatureBuf_657;
         Mult_Buf[69].Weight_n = Wgt_3_657;
         Mult_Buf[70].Feature_n = FeatureBuf_658;
         Mult_Buf[70].Weight_n = Wgt_3_658;
         Mult_Buf[71].Feature_n = FeatureBuf_659;
         Mult_Buf[71].Weight_n = Wgt_3_659;
         Mult_Buf[72].Feature_n = FeatureBuf_660;
         Mult_Buf[72].Weight_n = Wgt_3_660;
         Mult_Buf[73].Feature_n = FeatureBuf_661;
         Mult_Buf[73].Weight_n = Wgt_3_661;
         Mult_Buf[74].Feature_n = FeatureBuf_662;
         Mult_Buf[74].Weight_n = Wgt_3_662;
         Mult_Buf[75].Feature_n = FeatureBuf_663;
         Mult_Buf[75].Weight_n = Wgt_3_663;
         Mult_Buf[76].Feature_n = FeatureBuf_664;
         Mult_Buf[76].Weight_n = Wgt_3_664;
         Mult_Buf[77].Feature_n = FeatureBuf_665;
         Mult_Buf[77].Weight_n = Wgt_3_665;
         Mult_Buf[78].Feature_n = FeatureBuf_666;
         Mult_Buf[78].Weight_n = Wgt_3_666;
         Mult_Buf[79].Feature_n = FeatureBuf_667;
         Mult_Buf[79].Weight_n = Wgt_3_667;
         Mult_Buf[80].Feature_n = FeatureBuf_668;
         Mult_Buf[80].Weight_n = Wgt_3_668;
         Mult_Buf[81].Feature_n = FeatureBuf_669;
         Mult_Buf[81].Weight_n = Wgt_3_669;
         Mult_Buf[82].Feature_n = FeatureBuf_670;
         Mult_Buf[82].Weight_n = Wgt_3_670;
         Mult_Buf[83].Feature_n = FeatureBuf_671;
         Mult_Buf[83].Weight_n = Wgt_3_671;
         Mult_Buf[84].Feature_n = FeatureBuf_672;
         Mult_Buf[84].Weight_n = Wgt_3_672;
         Mult_Buf[85].Feature_n = FeatureBuf_673;
         Mult_Buf[85].Weight_n = Wgt_3_673;
         Mult_Buf[86].Feature_n = FeatureBuf_674;
         Mult_Buf[86].Weight_n = Wgt_3_674;
         Mult_Buf[87].Feature_n = FeatureBuf_675;
         Mult_Buf[87].Weight_n = Wgt_3_675;
         Mult_Buf[88].Feature_n = FeatureBuf_676;
         Mult_Buf[88].Weight_n = Wgt_3_676;
         Mult_Buf[89].Feature_n = FeatureBuf_677;
         Mult_Buf[89].Weight_n = Wgt_3_677;
         Mult_Buf[90].Feature_n = FeatureBuf_678;
         Mult_Buf[90].Weight_n = Wgt_3_678;
         Mult_Buf[91].Feature_n = FeatureBuf_679;
         Mult_Buf[91].Weight_n = Wgt_3_679;
         Mult_Buf[92].Feature_n = FeatureBuf_680;
         Mult_Buf[92].Weight_n = Wgt_3_680;
         Mult_Buf[93].Feature_n = FeatureBuf_681;
         Mult_Buf[93].Weight_n = Wgt_3_681;
         Mult_Buf[94].Feature_n = FeatureBuf_682;
         Mult_Buf[94].Weight_n = Wgt_3_682;
         Mult_Buf[95].Feature_n = FeatureBuf_683;
         Mult_Buf[95].Weight_n = Wgt_3_683;
         Mult_Buf[96].Feature_n = FeatureBuf_684;
         Mult_Buf[96].Weight_n = Wgt_3_684;
         Mult_Buf[97].Feature_n = FeatureBuf_685;
         Mult_Buf[97].Weight_n = Wgt_3_685;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     //Collect Partial result form Adder
         Res_1_0_n = Part_Res;
     end
    33:begin
     nxt_state = 34;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_686;
         Mult_Buf[0].Weight_n = Wgt_3_686;
         Mult_Buf[1].Feature_n = FeatureBuf_687;
         Mult_Buf[1].Weight_n = Wgt_3_687;
         Mult_Buf[2].Feature_n = FeatureBuf_688;
         Mult_Buf[2].Weight_n = Wgt_3_688;
         Mult_Buf[3].Feature_n = FeatureBuf_689;
         Mult_Buf[3].Weight_n = Wgt_3_689;
         Mult_Buf[4].Feature_n = FeatureBuf_690;
         Mult_Buf[4].Weight_n = Wgt_3_690;
         Mult_Buf[5].Feature_n = FeatureBuf_691;
         Mult_Buf[5].Weight_n = Wgt_3_691;
         Mult_Buf[6].Feature_n = FeatureBuf_692;
         Mult_Buf[6].Weight_n = Wgt_3_692;
         Mult_Buf[7].Feature_n = FeatureBuf_693;
         Mult_Buf[7].Weight_n = Wgt_3_693;
         Mult_Buf[8].Feature_n = FeatureBuf_694;
         Mult_Buf[8].Weight_n = Wgt_3_694;
         Mult_Buf[9].Feature_n = FeatureBuf_695;
         Mult_Buf[9].Weight_n = Wgt_3_695;
         Mult_Buf[10].Feature_n = FeatureBuf_696;
         Mult_Buf[10].Weight_n = Wgt_3_696;
         Mult_Buf[11].Feature_n = FeatureBuf_697;
         Mult_Buf[11].Weight_n = Wgt_3_697;
         Mult_Buf[12].Feature_n = FeatureBuf_698;
         Mult_Buf[12].Weight_n = Wgt_3_698;
         Mult_Buf[13].Feature_n = FeatureBuf_699;
         Mult_Buf[13].Weight_n = Wgt_3_699;
         Mult_Buf[14].Feature_n = FeatureBuf_700;
         Mult_Buf[14].Weight_n = Wgt_3_700;
         Mult_Buf[15].Feature_n = FeatureBuf_701;
         Mult_Buf[15].Weight_n = Wgt_3_701;
         Mult_Buf[16].Feature_n = FeatureBuf_702;
         Mult_Buf[16].Weight_n = Wgt_3_702;
         Mult_Buf[17].Feature_n = FeatureBuf_703;
         Mult_Buf[17].Weight_n = Wgt_3_703;
         Mult_Buf[18].Feature_n = FeatureBuf_704;
         Mult_Buf[18].Weight_n = Wgt_3_704;
         Mult_Buf[19].Feature_n = FeatureBuf_705;
         Mult_Buf[19].Weight_n = Wgt_3_705;
         Mult_Buf[20].Feature_n = FeatureBuf_706;
         Mult_Buf[20].Weight_n = Wgt_3_706;
         Mult_Buf[21].Feature_n = FeatureBuf_707;
         Mult_Buf[21].Weight_n = Wgt_3_707;
         Mult_Buf[22].Feature_n = FeatureBuf_708;
         Mult_Buf[22].Weight_n = Wgt_3_708;
         Mult_Buf[23].Feature_n = FeatureBuf_709;
         Mult_Buf[23].Weight_n = Wgt_3_709;
         Mult_Buf[24].Feature_n = FeatureBuf_710;
         Mult_Buf[24].Weight_n = Wgt_3_710;
         Mult_Buf[25].Feature_n = FeatureBuf_711;
         Mult_Buf[25].Weight_n = Wgt_3_711;
         Mult_Buf[26].Feature_n = FeatureBuf_712;
         Mult_Buf[26].Weight_n = Wgt_3_712;
         Mult_Buf[27].Feature_n = FeatureBuf_713;
         Mult_Buf[27].Weight_n = Wgt_3_713;
         Mult_Buf[28].Feature_n = FeatureBuf_714;
         Mult_Buf[28].Weight_n = Wgt_3_714;
         Mult_Buf[29].Feature_n = FeatureBuf_715;
         Mult_Buf[29].Weight_n = Wgt_3_715;
         Mult_Buf[30].Feature_n = FeatureBuf_716;
         Mult_Buf[30].Weight_n = Wgt_3_716;
         Mult_Buf[31].Feature_n = FeatureBuf_717;
         Mult_Buf[31].Weight_n = Wgt_3_717;
         Mult_Buf[32].Feature_n = FeatureBuf_718;
         Mult_Buf[32].Weight_n = Wgt_3_718;
         Mult_Buf[33].Feature_n = FeatureBuf_719;
         Mult_Buf[33].Weight_n = Wgt_3_719;
         Mult_Buf[34].Feature_n = FeatureBuf_720;
         Mult_Buf[34].Weight_n = Wgt_3_720;
         Mult_Buf[35].Feature_n = FeatureBuf_721;
         Mult_Buf[35].Weight_n = Wgt_3_721;
         Mult_Buf[36].Feature_n = FeatureBuf_722;
         Mult_Buf[36].Weight_n = Wgt_3_722;
         Mult_Buf[37].Feature_n = FeatureBuf_723;
         Mult_Buf[37].Weight_n = Wgt_3_723;
         Mult_Buf[38].Feature_n = FeatureBuf_724;
         Mult_Buf[38].Weight_n = Wgt_3_724;
         Mult_Buf[39].Feature_n = FeatureBuf_725;
         Mult_Buf[39].Weight_n = Wgt_3_725;
         Mult_Buf[40].Feature_n = FeatureBuf_726;
         Mult_Buf[40].Weight_n = Wgt_3_726;
         Mult_Buf[41].Feature_n = FeatureBuf_727;
         Mult_Buf[41].Weight_n = Wgt_3_727;
         Mult_Buf[42].Feature_n = FeatureBuf_728;
         Mult_Buf[42].Weight_n = Wgt_3_728;
         Mult_Buf[43].Feature_n = FeatureBuf_729;
         Mult_Buf[43].Weight_n = Wgt_3_729;
         Mult_Buf[44].Feature_n = FeatureBuf_730;
         Mult_Buf[44].Weight_n = Wgt_3_730;
         Mult_Buf[45].Feature_n = FeatureBuf_731;
         Mult_Buf[45].Weight_n = Wgt_3_731;
         Mult_Buf[46].Feature_n = FeatureBuf_732;
         Mult_Buf[46].Weight_n = Wgt_3_732;
         Mult_Buf[47].Feature_n = FeatureBuf_733;
         Mult_Buf[47].Weight_n = Wgt_3_733;
         Mult_Buf[48].Feature_n = FeatureBuf_734;
         Mult_Buf[48].Weight_n = Wgt_3_734;
         Mult_Buf[49].Feature_n = FeatureBuf_735;
         Mult_Buf[49].Weight_n = Wgt_3_735;
         Mult_Buf[50].Feature_n = FeatureBuf_736;
         Mult_Buf[50].Weight_n = Wgt_3_736;
         Mult_Buf[51].Feature_n = FeatureBuf_737;
         Mult_Buf[51].Weight_n = Wgt_3_737;
         Mult_Buf[52].Feature_n = FeatureBuf_738;
         Mult_Buf[52].Weight_n = Wgt_3_738;
         Mult_Buf[53].Feature_n = FeatureBuf_739;
         Mult_Buf[53].Weight_n = Wgt_3_739;
         Mult_Buf[54].Feature_n = FeatureBuf_740;
         Mult_Buf[54].Weight_n = Wgt_3_740;
         Mult_Buf[55].Feature_n = FeatureBuf_741;
         Mult_Buf[55].Weight_n = Wgt_3_741;
         Mult_Buf[56].Feature_n = FeatureBuf_742;
         Mult_Buf[56].Weight_n = Wgt_3_742;
         Mult_Buf[57].Feature_n = FeatureBuf_743;
         Mult_Buf[57].Weight_n = Wgt_3_743;
         Mult_Buf[58].Feature_n = FeatureBuf_744;
         Mult_Buf[58].Weight_n = Wgt_3_744;
         Mult_Buf[59].Feature_n = FeatureBuf_745;
         Mult_Buf[59].Weight_n = Wgt_3_745;
         Mult_Buf[60].Feature_n = FeatureBuf_746;
         Mult_Buf[60].Weight_n = Wgt_3_746;
         Mult_Buf[61].Feature_n = FeatureBuf_747;
         Mult_Buf[61].Weight_n = Wgt_3_747;
         Mult_Buf[62].Feature_n = FeatureBuf_748;
         Mult_Buf[62].Weight_n = Wgt_3_748;
         Mult_Buf[63].Feature_n = FeatureBuf_749;
         Mult_Buf[63].Weight_n = Wgt_3_749;
         Mult_Buf[64].Feature_n = FeatureBuf_750;
         Mult_Buf[64].Weight_n = Wgt_3_750;
         Mult_Buf[65].Feature_n = FeatureBuf_751;
         Mult_Buf[65].Weight_n = Wgt_3_751;
         Mult_Buf[66].Feature_n = FeatureBuf_752;
         Mult_Buf[66].Weight_n = Wgt_3_752;
         Mult_Buf[67].Feature_n = FeatureBuf_753;
         Mult_Buf[67].Weight_n = Wgt_3_753;
         Mult_Buf[68].Feature_n = FeatureBuf_754;
         Mult_Buf[68].Weight_n = Wgt_3_754;
         Mult_Buf[69].Feature_n = FeatureBuf_755;
         Mult_Buf[69].Weight_n = Wgt_3_755;
         Mult_Buf[70].Feature_n = FeatureBuf_756;
         Mult_Buf[70].Weight_n = Wgt_3_756;
         Mult_Buf[71].Feature_n = FeatureBuf_757;
         Mult_Buf[71].Weight_n = Wgt_3_757;
         Mult_Buf[72].Feature_n = FeatureBuf_758;
         Mult_Buf[72].Weight_n = Wgt_3_758;
         Mult_Buf[73].Feature_n = FeatureBuf_759;
         Mult_Buf[73].Weight_n = Wgt_3_759;
         Mult_Buf[74].Feature_n = FeatureBuf_760;
         Mult_Buf[74].Weight_n = Wgt_3_760;
         Mult_Buf[75].Feature_n = FeatureBuf_761;
         Mult_Buf[75].Weight_n = Wgt_3_761;
         Mult_Buf[76].Feature_n = FeatureBuf_762;
         Mult_Buf[76].Weight_n = Wgt_3_762;
         Mult_Buf[77].Feature_n = FeatureBuf_763;
         Mult_Buf[77].Weight_n = Wgt_3_763;
         Mult_Buf[78].Feature_n = FeatureBuf_764;
         Mult_Buf[78].Weight_n = Wgt_3_764;
         Mult_Buf[79].Feature_n = FeatureBuf_765;
         Mult_Buf[79].Weight_n = Wgt_3_765;
         Mult_Buf[80].Feature_n = FeatureBuf_766;
         Mult_Buf[80].Weight_n = Wgt_3_766;
         Mult_Buf[81].Feature_n = FeatureBuf_767;
         Mult_Buf[81].Weight_n = Wgt_3_767;
         Mult_Buf[82].Feature_n = FeatureBuf_768;
         Mult_Buf[82].Weight_n = Wgt_3_768;
         Mult_Buf[83].Feature_n = FeatureBuf_769;
         Mult_Buf[83].Weight_n = Wgt_3_769;
         Mult_Buf[84].Feature_n = FeatureBuf_770;
         Mult_Buf[84].Weight_n = Wgt_3_770;
         Mult_Buf[85].Feature_n = FeatureBuf_771;
         Mult_Buf[85].Weight_n = Wgt_3_771;
         Mult_Buf[86].Feature_n = FeatureBuf_772;
         Mult_Buf[86].Weight_n = Wgt_3_772;
         Mult_Buf[87].Feature_n = FeatureBuf_773;
         Mult_Buf[87].Weight_n = Wgt_3_773;
         Mult_Buf[88].Feature_n = FeatureBuf_774;
         Mult_Buf[88].Weight_n = Wgt_3_774;
         Mult_Buf[89].Feature_n = FeatureBuf_775;
         Mult_Buf[89].Weight_n = Wgt_3_775;
         Mult_Buf[90].Feature_n = FeatureBuf_776;
         Mult_Buf[90].Weight_n = Wgt_3_776;
         Mult_Buf[91].Feature_n = FeatureBuf_777;
         Mult_Buf[91].Weight_n = Wgt_3_777;
         Mult_Buf[92].Feature_n = FeatureBuf_778;
         Mult_Buf[92].Weight_n = Wgt_3_778;
         Mult_Buf[93].Feature_n = FeatureBuf_779;
         Mult_Buf[93].Weight_n = Wgt_3_779;
         Mult_Buf[94].Feature_n = FeatureBuf_780;
         Mult_Buf[94].Weight_n = Wgt_3_780;
         Mult_Buf[95].Feature_n = FeatureBuf_781;
         Mult_Buf[95].Weight_n = Wgt_3_781;
         Mult_Buf[96].Feature_n = FeatureBuf_782;
         Mult_Buf[96].Weight_n = Wgt_3_782;
         Mult_Buf[97].Feature_n = FeatureBuf_783;
         Mult_Buf[97].Weight_n = Wgt_3_783;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     //Collect Partial result form Adder
         Res_1_1_n = Part_Res;
     end
    34:begin
     nxt_state = 35;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_0;
         Mult_Buf[0].Weight_n = Wgt_4_0;
         Mult_Buf[1].Feature_n = FeatureBuf_1;
         Mult_Buf[1].Weight_n = Wgt_4_1;
         Mult_Buf[2].Feature_n = FeatureBuf_2;
         Mult_Buf[2].Weight_n = Wgt_4_2;
         Mult_Buf[3].Feature_n = FeatureBuf_3;
         Mult_Buf[3].Weight_n = Wgt_4_3;
         Mult_Buf[4].Feature_n = FeatureBuf_4;
         Mult_Buf[4].Weight_n = Wgt_4_4;
         Mult_Buf[5].Feature_n = FeatureBuf_5;
         Mult_Buf[5].Weight_n = Wgt_4_5;
         Mult_Buf[6].Feature_n = FeatureBuf_6;
         Mult_Buf[6].Weight_n = Wgt_4_6;
         Mult_Buf[7].Feature_n = FeatureBuf_7;
         Mult_Buf[7].Weight_n = Wgt_4_7;
         Mult_Buf[8].Feature_n = FeatureBuf_8;
         Mult_Buf[8].Weight_n = Wgt_4_8;
         Mult_Buf[9].Feature_n = FeatureBuf_9;
         Mult_Buf[9].Weight_n = Wgt_4_9;
         Mult_Buf[10].Feature_n = FeatureBuf_10;
         Mult_Buf[10].Weight_n = Wgt_4_10;
         Mult_Buf[11].Feature_n = FeatureBuf_11;
         Mult_Buf[11].Weight_n = Wgt_4_11;
         Mult_Buf[12].Feature_n = FeatureBuf_12;
         Mult_Buf[12].Weight_n = Wgt_4_12;
         Mult_Buf[13].Feature_n = FeatureBuf_13;
         Mult_Buf[13].Weight_n = Wgt_4_13;
         Mult_Buf[14].Feature_n = FeatureBuf_14;
         Mult_Buf[14].Weight_n = Wgt_4_14;
         Mult_Buf[15].Feature_n = FeatureBuf_15;
         Mult_Buf[15].Weight_n = Wgt_4_15;
         Mult_Buf[16].Feature_n = FeatureBuf_16;
         Mult_Buf[16].Weight_n = Wgt_4_16;
         Mult_Buf[17].Feature_n = FeatureBuf_17;
         Mult_Buf[17].Weight_n = Wgt_4_17;
         Mult_Buf[18].Feature_n = FeatureBuf_18;
         Mult_Buf[18].Weight_n = Wgt_4_18;
         Mult_Buf[19].Feature_n = FeatureBuf_19;
         Mult_Buf[19].Weight_n = Wgt_4_19;
         Mult_Buf[20].Feature_n = FeatureBuf_20;
         Mult_Buf[20].Weight_n = Wgt_4_20;
         Mult_Buf[21].Feature_n = FeatureBuf_21;
         Mult_Buf[21].Weight_n = Wgt_4_21;
         Mult_Buf[22].Feature_n = FeatureBuf_22;
         Mult_Buf[22].Weight_n = Wgt_4_22;
         Mult_Buf[23].Feature_n = FeatureBuf_23;
         Mult_Buf[23].Weight_n = Wgt_4_23;
         Mult_Buf[24].Feature_n = FeatureBuf_24;
         Mult_Buf[24].Weight_n = Wgt_4_24;
         Mult_Buf[25].Feature_n = FeatureBuf_25;
         Mult_Buf[25].Weight_n = Wgt_4_25;
         Mult_Buf[26].Feature_n = FeatureBuf_26;
         Mult_Buf[26].Weight_n = Wgt_4_26;
         Mult_Buf[27].Feature_n = FeatureBuf_27;
         Mult_Buf[27].Weight_n = Wgt_4_27;
         Mult_Buf[28].Feature_n = FeatureBuf_28;
         Mult_Buf[28].Weight_n = Wgt_4_28;
         Mult_Buf[29].Feature_n = FeatureBuf_29;
         Mult_Buf[29].Weight_n = Wgt_4_29;
         Mult_Buf[30].Feature_n = FeatureBuf_30;
         Mult_Buf[30].Weight_n = Wgt_4_30;
         Mult_Buf[31].Feature_n = FeatureBuf_31;
         Mult_Buf[31].Weight_n = Wgt_4_31;
         Mult_Buf[32].Feature_n = FeatureBuf_32;
         Mult_Buf[32].Weight_n = Wgt_4_32;
         Mult_Buf[33].Feature_n = FeatureBuf_33;
         Mult_Buf[33].Weight_n = Wgt_4_33;
         Mult_Buf[34].Feature_n = FeatureBuf_34;
         Mult_Buf[34].Weight_n = Wgt_4_34;
         Mult_Buf[35].Feature_n = FeatureBuf_35;
         Mult_Buf[35].Weight_n = Wgt_4_35;
         Mult_Buf[36].Feature_n = FeatureBuf_36;
         Mult_Buf[36].Weight_n = Wgt_4_36;
         Mult_Buf[37].Feature_n = FeatureBuf_37;
         Mult_Buf[37].Weight_n = Wgt_4_37;
         Mult_Buf[38].Feature_n = FeatureBuf_38;
         Mult_Buf[38].Weight_n = Wgt_4_38;
         Mult_Buf[39].Feature_n = FeatureBuf_39;
         Mult_Buf[39].Weight_n = Wgt_4_39;
         Mult_Buf[40].Feature_n = FeatureBuf_40;
         Mult_Buf[40].Weight_n = Wgt_4_40;
         Mult_Buf[41].Feature_n = FeatureBuf_41;
         Mult_Buf[41].Weight_n = Wgt_4_41;
         Mult_Buf[42].Feature_n = FeatureBuf_42;
         Mult_Buf[42].Weight_n = Wgt_4_42;
         Mult_Buf[43].Feature_n = FeatureBuf_43;
         Mult_Buf[43].Weight_n = Wgt_4_43;
         Mult_Buf[44].Feature_n = FeatureBuf_44;
         Mult_Buf[44].Weight_n = Wgt_4_44;
         Mult_Buf[45].Feature_n = FeatureBuf_45;
         Mult_Buf[45].Weight_n = Wgt_4_45;
         Mult_Buf[46].Feature_n = FeatureBuf_46;
         Mult_Buf[46].Weight_n = Wgt_4_46;
         Mult_Buf[47].Feature_n = FeatureBuf_47;
         Mult_Buf[47].Weight_n = Wgt_4_47;
         Mult_Buf[48].Feature_n = FeatureBuf_48;
         Mult_Buf[48].Weight_n = Wgt_4_48;
         Mult_Buf[49].Feature_n = FeatureBuf_49;
         Mult_Buf[49].Weight_n = Wgt_4_49;
         Mult_Buf[50].Feature_n = FeatureBuf_50;
         Mult_Buf[50].Weight_n = Wgt_4_50;
         Mult_Buf[51].Feature_n = FeatureBuf_51;
         Mult_Buf[51].Weight_n = Wgt_4_51;
         Mult_Buf[52].Feature_n = FeatureBuf_52;
         Mult_Buf[52].Weight_n = Wgt_4_52;
         Mult_Buf[53].Feature_n = FeatureBuf_53;
         Mult_Buf[53].Weight_n = Wgt_4_53;
         Mult_Buf[54].Feature_n = FeatureBuf_54;
         Mult_Buf[54].Weight_n = Wgt_4_54;
         Mult_Buf[55].Feature_n = FeatureBuf_55;
         Mult_Buf[55].Weight_n = Wgt_4_55;
         Mult_Buf[56].Feature_n = FeatureBuf_56;
         Mult_Buf[56].Weight_n = Wgt_4_56;
         Mult_Buf[57].Feature_n = FeatureBuf_57;
         Mult_Buf[57].Weight_n = Wgt_4_57;
         Mult_Buf[58].Feature_n = FeatureBuf_58;
         Mult_Buf[58].Weight_n = Wgt_4_58;
         Mult_Buf[59].Feature_n = FeatureBuf_59;
         Mult_Buf[59].Weight_n = Wgt_4_59;
         Mult_Buf[60].Feature_n = FeatureBuf_60;
         Mult_Buf[60].Weight_n = Wgt_4_60;
         Mult_Buf[61].Feature_n = FeatureBuf_61;
         Mult_Buf[61].Weight_n = Wgt_4_61;
         Mult_Buf[62].Feature_n = FeatureBuf_62;
         Mult_Buf[62].Weight_n = Wgt_4_62;
         Mult_Buf[63].Feature_n = FeatureBuf_63;
         Mult_Buf[63].Weight_n = Wgt_4_63;
         Mult_Buf[64].Feature_n = FeatureBuf_64;
         Mult_Buf[64].Weight_n = Wgt_4_64;
         Mult_Buf[65].Feature_n = FeatureBuf_65;
         Mult_Buf[65].Weight_n = Wgt_4_65;
         Mult_Buf[66].Feature_n = FeatureBuf_66;
         Mult_Buf[66].Weight_n = Wgt_4_66;
         Mult_Buf[67].Feature_n = FeatureBuf_67;
         Mult_Buf[67].Weight_n = Wgt_4_67;
         Mult_Buf[68].Feature_n = FeatureBuf_68;
         Mult_Buf[68].Weight_n = Wgt_4_68;
         Mult_Buf[69].Feature_n = FeatureBuf_69;
         Mult_Buf[69].Weight_n = Wgt_4_69;
         Mult_Buf[70].Feature_n = FeatureBuf_70;
         Mult_Buf[70].Weight_n = Wgt_4_70;
         Mult_Buf[71].Feature_n = FeatureBuf_71;
         Mult_Buf[71].Weight_n = Wgt_4_71;
         Mult_Buf[72].Feature_n = FeatureBuf_72;
         Mult_Buf[72].Weight_n = Wgt_4_72;
         Mult_Buf[73].Feature_n = FeatureBuf_73;
         Mult_Buf[73].Weight_n = Wgt_4_73;
         Mult_Buf[74].Feature_n = FeatureBuf_74;
         Mult_Buf[74].Weight_n = Wgt_4_74;
         Mult_Buf[75].Feature_n = FeatureBuf_75;
         Mult_Buf[75].Weight_n = Wgt_4_75;
         Mult_Buf[76].Feature_n = FeatureBuf_76;
         Mult_Buf[76].Weight_n = Wgt_4_76;
         Mult_Buf[77].Feature_n = FeatureBuf_77;
         Mult_Buf[77].Weight_n = Wgt_4_77;
         Mult_Buf[78].Feature_n = FeatureBuf_78;
         Mult_Buf[78].Weight_n = Wgt_4_78;
         Mult_Buf[79].Feature_n = FeatureBuf_79;
         Mult_Buf[79].Weight_n = Wgt_4_79;
         Mult_Buf[80].Feature_n = FeatureBuf_80;
         Mult_Buf[80].Weight_n = Wgt_4_80;
         Mult_Buf[81].Feature_n = FeatureBuf_81;
         Mult_Buf[81].Weight_n = Wgt_4_81;
         Mult_Buf[82].Feature_n = FeatureBuf_82;
         Mult_Buf[82].Weight_n = Wgt_4_82;
         Mult_Buf[83].Feature_n = FeatureBuf_83;
         Mult_Buf[83].Weight_n = Wgt_4_83;
         Mult_Buf[84].Feature_n = FeatureBuf_84;
         Mult_Buf[84].Weight_n = Wgt_4_84;
         Mult_Buf[85].Feature_n = FeatureBuf_85;
         Mult_Buf[85].Weight_n = Wgt_4_85;
         Mult_Buf[86].Feature_n = FeatureBuf_86;
         Mult_Buf[86].Weight_n = Wgt_4_86;
         Mult_Buf[87].Feature_n = FeatureBuf_87;
         Mult_Buf[87].Weight_n = Wgt_4_87;
         Mult_Buf[88].Feature_n = FeatureBuf_88;
         Mult_Buf[88].Weight_n = Wgt_4_88;
         Mult_Buf[89].Feature_n = FeatureBuf_89;
         Mult_Buf[89].Weight_n = Wgt_4_89;
         Mult_Buf[90].Feature_n = FeatureBuf_90;
         Mult_Buf[90].Weight_n = Wgt_4_90;
         Mult_Buf[91].Feature_n = FeatureBuf_91;
         Mult_Buf[91].Weight_n = Wgt_4_91;
         Mult_Buf[92].Feature_n = FeatureBuf_92;
         Mult_Buf[92].Weight_n = Wgt_4_92;
         Mult_Buf[93].Feature_n = FeatureBuf_93;
         Mult_Buf[93].Weight_n = Wgt_4_93;
         Mult_Buf[94].Feature_n = FeatureBuf_94;
         Mult_Buf[94].Weight_n = Wgt_4_94;
         Mult_Buf[95].Feature_n = FeatureBuf_95;
         Mult_Buf[95].Weight_n = Wgt_4_95;
         Mult_Buf[96].Feature_n = FeatureBuf_96;
         Mult_Buf[96].Weight_n = Wgt_4_96;
         Mult_Buf[97].Feature_n = FeatureBuf_97;
         Mult_Buf[97].Weight_n = Wgt_4_97;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     //Collect Partial result form Adder
         Res_1_2_n = Part_Res;
     end
    35:begin
     nxt_state = 36;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_98;
         Mult_Buf[0].Weight_n = Wgt_4_98;
         Mult_Buf[1].Feature_n = FeatureBuf_99;
         Mult_Buf[1].Weight_n = Wgt_4_99;
         Mult_Buf[2].Feature_n = FeatureBuf_100;
         Mult_Buf[2].Weight_n = Wgt_4_100;
         Mult_Buf[3].Feature_n = FeatureBuf_101;
         Mult_Buf[3].Weight_n = Wgt_4_101;
         Mult_Buf[4].Feature_n = FeatureBuf_102;
         Mult_Buf[4].Weight_n = Wgt_4_102;
         Mult_Buf[5].Feature_n = FeatureBuf_103;
         Mult_Buf[5].Weight_n = Wgt_4_103;
         Mult_Buf[6].Feature_n = FeatureBuf_104;
         Mult_Buf[6].Weight_n = Wgt_4_104;
         Mult_Buf[7].Feature_n = FeatureBuf_105;
         Mult_Buf[7].Weight_n = Wgt_4_105;
         Mult_Buf[8].Feature_n = FeatureBuf_106;
         Mult_Buf[8].Weight_n = Wgt_4_106;
         Mult_Buf[9].Feature_n = FeatureBuf_107;
         Mult_Buf[9].Weight_n = Wgt_4_107;
         Mult_Buf[10].Feature_n = FeatureBuf_108;
         Mult_Buf[10].Weight_n = Wgt_4_108;
         Mult_Buf[11].Feature_n = FeatureBuf_109;
         Mult_Buf[11].Weight_n = Wgt_4_109;
         Mult_Buf[12].Feature_n = FeatureBuf_110;
         Mult_Buf[12].Weight_n = Wgt_4_110;
         Mult_Buf[13].Feature_n = FeatureBuf_111;
         Mult_Buf[13].Weight_n = Wgt_4_111;
         Mult_Buf[14].Feature_n = FeatureBuf_112;
         Mult_Buf[14].Weight_n = Wgt_4_112;
         Mult_Buf[15].Feature_n = FeatureBuf_113;
         Mult_Buf[15].Weight_n = Wgt_4_113;
         Mult_Buf[16].Feature_n = FeatureBuf_114;
         Mult_Buf[16].Weight_n = Wgt_4_114;
         Mult_Buf[17].Feature_n = FeatureBuf_115;
         Mult_Buf[17].Weight_n = Wgt_4_115;
         Mult_Buf[18].Feature_n = FeatureBuf_116;
         Mult_Buf[18].Weight_n = Wgt_4_116;
         Mult_Buf[19].Feature_n = FeatureBuf_117;
         Mult_Buf[19].Weight_n = Wgt_4_117;
         Mult_Buf[20].Feature_n = FeatureBuf_118;
         Mult_Buf[20].Weight_n = Wgt_4_118;
         Mult_Buf[21].Feature_n = FeatureBuf_119;
         Mult_Buf[21].Weight_n = Wgt_4_119;
         Mult_Buf[22].Feature_n = FeatureBuf_120;
         Mult_Buf[22].Weight_n = Wgt_4_120;
         Mult_Buf[23].Feature_n = FeatureBuf_121;
         Mult_Buf[23].Weight_n = Wgt_4_121;
         Mult_Buf[24].Feature_n = FeatureBuf_122;
         Mult_Buf[24].Weight_n = Wgt_4_122;
         Mult_Buf[25].Feature_n = FeatureBuf_123;
         Mult_Buf[25].Weight_n = Wgt_4_123;
         Mult_Buf[26].Feature_n = FeatureBuf_124;
         Mult_Buf[26].Weight_n = Wgt_4_124;
         Mult_Buf[27].Feature_n = FeatureBuf_125;
         Mult_Buf[27].Weight_n = Wgt_4_125;
         Mult_Buf[28].Feature_n = FeatureBuf_126;
         Mult_Buf[28].Weight_n = Wgt_4_126;
         Mult_Buf[29].Feature_n = FeatureBuf_127;
         Mult_Buf[29].Weight_n = Wgt_4_127;
         Mult_Buf[30].Feature_n = FeatureBuf_128;
         Mult_Buf[30].Weight_n = Wgt_4_128;
         Mult_Buf[31].Feature_n = FeatureBuf_129;
         Mult_Buf[31].Weight_n = Wgt_4_129;
         Mult_Buf[32].Feature_n = FeatureBuf_130;
         Mult_Buf[32].Weight_n = Wgt_4_130;
         Mult_Buf[33].Feature_n = FeatureBuf_131;
         Mult_Buf[33].Weight_n = Wgt_4_131;
         Mult_Buf[34].Feature_n = FeatureBuf_132;
         Mult_Buf[34].Weight_n = Wgt_4_132;
         Mult_Buf[35].Feature_n = FeatureBuf_133;
         Mult_Buf[35].Weight_n = Wgt_4_133;
         Mult_Buf[36].Feature_n = FeatureBuf_134;
         Mult_Buf[36].Weight_n = Wgt_4_134;
         Mult_Buf[37].Feature_n = FeatureBuf_135;
         Mult_Buf[37].Weight_n = Wgt_4_135;
         Mult_Buf[38].Feature_n = FeatureBuf_136;
         Mult_Buf[38].Weight_n = Wgt_4_136;
         Mult_Buf[39].Feature_n = FeatureBuf_137;
         Mult_Buf[39].Weight_n = Wgt_4_137;
         Mult_Buf[40].Feature_n = FeatureBuf_138;
         Mult_Buf[40].Weight_n = Wgt_4_138;
         Mult_Buf[41].Feature_n = FeatureBuf_139;
         Mult_Buf[41].Weight_n = Wgt_4_139;
         Mult_Buf[42].Feature_n = FeatureBuf_140;
         Mult_Buf[42].Weight_n = Wgt_4_140;
         Mult_Buf[43].Feature_n = FeatureBuf_141;
         Mult_Buf[43].Weight_n = Wgt_4_141;
         Mult_Buf[44].Feature_n = FeatureBuf_142;
         Mult_Buf[44].Weight_n = Wgt_4_142;
         Mult_Buf[45].Feature_n = FeatureBuf_143;
         Mult_Buf[45].Weight_n = Wgt_4_143;
         Mult_Buf[46].Feature_n = FeatureBuf_144;
         Mult_Buf[46].Weight_n = Wgt_4_144;
         Mult_Buf[47].Feature_n = FeatureBuf_145;
         Mult_Buf[47].Weight_n = Wgt_4_145;
         Mult_Buf[48].Feature_n = FeatureBuf_146;
         Mult_Buf[48].Weight_n = Wgt_4_146;
         Mult_Buf[49].Feature_n = FeatureBuf_147;
         Mult_Buf[49].Weight_n = Wgt_4_147;
         Mult_Buf[50].Feature_n = FeatureBuf_148;
         Mult_Buf[50].Weight_n = Wgt_4_148;
         Mult_Buf[51].Feature_n = FeatureBuf_149;
         Mult_Buf[51].Weight_n = Wgt_4_149;
         Mult_Buf[52].Feature_n = FeatureBuf_150;
         Mult_Buf[52].Weight_n = Wgt_4_150;
         Mult_Buf[53].Feature_n = FeatureBuf_151;
         Mult_Buf[53].Weight_n = Wgt_4_151;
         Mult_Buf[54].Feature_n = FeatureBuf_152;
         Mult_Buf[54].Weight_n = Wgt_4_152;
         Mult_Buf[55].Feature_n = FeatureBuf_153;
         Mult_Buf[55].Weight_n = Wgt_4_153;
         Mult_Buf[56].Feature_n = FeatureBuf_154;
         Mult_Buf[56].Weight_n = Wgt_4_154;
         Mult_Buf[57].Feature_n = FeatureBuf_155;
         Mult_Buf[57].Weight_n = Wgt_4_155;
         Mult_Buf[58].Feature_n = FeatureBuf_156;
         Mult_Buf[58].Weight_n = Wgt_4_156;
         Mult_Buf[59].Feature_n = FeatureBuf_157;
         Mult_Buf[59].Weight_n = Wgt_4_157;
         Mult_Buf[60].Feature_n = FeatureBuf_158;
         Mult_Buf[60].Weight_n = Wgt_4_158;
         Mult_Buf[61].Feature_n = FeatureBuf_159;
         Mult_Buf[61].Weight_n = Wgt_4_159;
         Mult_Buf[62].Feature_n = FeatureBuf_160;
         Mult_Buf[62].Weight_n = Wgt_4_160;
         Mult_Buf[63].Feature_n = FeatureBuf_161;
         Mult_Buf[63].Weight_n = Wgt_4_161;
         Mult_Buf[64].Feature_n = FeatureBuf_162;
         Mult_Buf[64].Weight_n = Wgt_4_162;
         Mult_Buf[65].Feature_n = FeatureBuf_163;
         Mult_Buf[65].Weight_n = Wgt_4_163;
         Mult_Buf[66].Feature_n = FeatureBuf_164;
         Mult_Buf[66].Weight_n = Wgt_4_164;
         Mult_Buf[67].Feature_n = FeatureBuf_165;
         Mult_Buf[67].Weight_n = Wgt_4_165;
         Mult_Buf[68].Feature_n = FeatureBuf_166;
         Mult_Buf[68].Weight_n = Wgt_4_166;
         Mult_Buf[69].Feature_n = FeatureBuf_167;
         Mult_Buf[69].Weight_n = Wgt_4_167;
         Mult_Buf[70].Feature_n = FeatureBuf_168;
         Mult_Buf[70].Weight_n = Wgt_4_168;
         Mult_Buf[71].Feature_n = FeatureBuf_169;
         Mult_Buf[71].Weight_n = Wgt_4_169;
         Mult_Buf[72].Feature_n = FeatureBuf_170;
         Mult_Buf[72].Weight_n = Wgt_4_170;
         Mult_Buf[73].Feature_n = FeatureBuf_171;
         Mult_Buf[73].Weight_n = Wgt_4_171;
         Mult_Buf[74].Feature_n = FeatureBuf_172;
         Mult_Buf[74].Weight_n = Wgt_4_172;
         Mult_Buf[75].Feature_n = FeatureBuf_173;
         Mult_Buf[75].Weight_n = Wgt_4_173;
         Mult_Buf[76].Feature_n = FeatureBuf_174;
         Mult_Buf[76].Weight_n = Wgt_4_174;
         Mult_Buf[77].Feature_n = FeatureBuf_175;
         Mult_Buf[77].Weight_n = Wgt_4_175;
         Mult_Buf[78].Feature_n = FeatureBuf_176;
         Mult_Buf[78].Weight_n = Wgt_4_176;
         Mult_Buf[79].Feature_n = FeatureBuf_177;
         Mult_Buf[79].Weight_n = Wgt_4_177;
         Mult_Buf[80].Feature_n = FeatureBuf_178;
         Mult_Buf[80].Weight_n = Wgt_4_178;
         Mult_Buf[81].Feature_n = FeatureBuf_179;
         Mult_Buf[81].Weight_n = Wgt_4_179;
         Mult_Buf[82].Feature_n = FeatureBuf_180;
         Mult_Buf[82].Weight_n = Wgt_4_180;
         Mult_Buf[83].Feature_n = FeatureBuf_181;
         Mult_Buf[83].Weight_n = Wgt_4_181;
         Mult_Buf[84].Feature_n = FeatureBuf_182;
         Mult_Buf[84].Weight_n = Wgt_4_182;
         Mult_Buf[85].Feature_n = FeatureBuf_183;
         Mult_Buf[85].Weight_n = Wgt_4_183;
         Mult_Buf[86].Feature_n = FeatureBuf_184;
         Mult_Buf[86].Weight_n = Wgt_4_184;
         Mult_Buf[87].Feature_n = FeatureBuf_185;
         Mult_Buf[87].Weight_n = Wgt_4_185;
         Mult_Buf[88].Feature_n = FeatureBuf_186;
         Mult_Buf[88].Weight_n = Wgt_4_186;
         Mult_Buf[89].Feature_n = FeatureBuf_187;
         Mult_Buf[89].Weight_n = Wgt_4_187;
         Mult_Buf[90].Feature_n = FeatureBuf_188;
         Mult_Buf[90].Weight_n = Wgt_4_188;
         Mult_Buf[91].Feature_n = FeatureBuf_189;
         Mult_Buf[91].Weight_n = Wgt_4_189;
         Mult_Buf[92].Feature_n = FeatureBuf_190;
         Mult_Buf[92].Weight_n = Wgt_4_190;
         Mult_Buf[93].Feature_n = FeatureBuf_191;
         Mult_Buf[93].Weight_n = Wgt_4_191;
         Mult_Buf[94].Feature_n = FeatureBuf_192;
         Mult_Buf[94].Weight_n = Wgt_4_192;
         Mult_Buf[95].Feature_n = FeatureBuf_193;
         Mult_Buf[95].Weight_n = Wgt_4_193;
         Mult_Buf[96].Feature_n = FeatureBuf_194;
         Mult_Buf[96].Weight_n = Wgt_4_194;
         Mult_Buf[97].Feature_n = FeatureBuf_195;
         Mult_Buf[97].Weight_n = Wgt_4_195;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     //Collect Partial result form Adder
         Res_1_3_n = Part_Res;
     end
    36:begin
     nxt_state = 37;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_196;
         Mult_Buf[0].Weight_n = Wgt_4_196;
         Mult_Buf[1].Feature_n = FeatureBuf_197;
         Mult_Buf[1].Weight_n = Wgt_4_197;
         Mult_Buf[2].Feature_n = FeatureBuf_198;
         Mult_Buf[2].Weight_n = Wgt_4_198;
         Mult_Buf[3].Feature_n = FeatureBuf_199;
         Mult_Buf[3].Weight_n = Wgt_4_199;
         Mult_Buf[4].Feature_n = FeatureBuf_200;
         Mult_Buf[4].Weight_n = Wgt_4_200;
         Mult_Buf[5].Feature_n = FeatureBuf_201;
         Mult_Buf[5].Weight_n = Wgt_4_201;
         Mult_Buf[6].Feature_n = FeatureBuf_202;
         Mult_Buf[6].Weight_n = Wgt_4_202;
         Mult_Buf[7].Feature_n = FeatureBuf_203;
         Mult_Buf[7].Weight_n = Wgt_4_203;
         Mult_Buf[8].Feature_n = FeatureBuf_204;
         Mult_Buf[8].Weight_n = Wgt_4_204;
         Mult_Buf[9].Feature_n = FeatureBuf_205;
         Mult_Buf[9].Weight_n = Wgt_4_205;
         Mult_Buf[10].Feature_n = FeatureBuf_206;
         Mult_Buf[10].Weight_n = Wgt_4_206;
         Mult_Buf[11].Feature_n = FeatureBuf_207;
         Mult_Buf[11].Weight_n = Wgt_4_207;
         Mult_Buf[12].Feature_n = FeatureBuf_208;
         Mult_Buf[12].Weight_n = Wgt_4_208;
         Mult_Buf[13].Feature_n = FeatureBuf_209;
         Mult_Buf[13].Weight_n = Wgt_4_209;
         Mult_Buf[14].Feature_n = FeatureBuf_210;
         Mult_Buf[14].Weight_n = Wgt_4_210;
         Mult_Buf[15].Feature_n = FeatureBuf_211;
         Mult_Buf[15].Weight_n = Wgt_4_211;
         Mult_Buf[16].Feature_n = FeatureBuf_212;
         Mult_Buf[16].Weight_n = Wgt_4_212;
         Mult_Buf[17].Feature_n = FeatureBuf_213;
         Mult_Buf[17].Weight_n = Wgt_4_213;
         Mult_Buf[18].Feature_n = FeatureBuf_214;
         Mult_Buf[18].Weight_n = Wgt_4_214;
         Mult_Buf[19].Feature_n = FeatureBuf_215;
         Mult_Buf[19].Weight_n = Wgt_4_215;
         Mult_Buf[20].Feature_n = FeatureBuf_216;
         Mult_Buf[20].Weight_n = Wgt_4_216;
         Mult_Buf[21].Feature_n = FeatureBuf_217;
         Mult_Buf[21].Weight_n = Wgt_4_217;
         Mult_Buf[22].Feature_n = FeatureBuf_218;
         Mult_Buf[22].Weight_n = Wgt_4_218;
         Mult_Buf[23].Feature_n = FeatureBuf_219;
         Mult_Buf[23].Weight_n = Wgt_4_219;
         Mult_Buf[24].Feature_n = FeatureBuf_220;
         Mult_Buf[24].Weight_n = Wgt_4_220;
         Mult_Buf[25].Feature_n = FeatureBuf_221;
         Mult_Buf[25].Weight_n = Wgt_4_221;
         Mult_Buf[26].Feature_n = FeatureBuf_222;
         Mult_Buf[26].Weight_n = Wgt_4_222;
         Mult_Buf[27].Feature_n = FeatureBuf_223;
         Mult_Buf[27].Weight_n = Wgt_4_223;
         Mult_Buf[28].Feature_n = FeatureBuf_224;
         Mult_Buf[28].Weight_n = Wgt_4_224;
         Mult_Buf[29].Feature_n = FeatureBuf_225;
         Mult_Buf[29].Weight_n = Wgt_4_225;
         Mult_Buf[30].Feature_n = FeatureBuf_226;
         Mult_Buf[30].Weight_n = Wgt_4_226;
         Mult_Buf[31].Feature_n = FeatureBuf_227;
         Mult_Buf[31].Weight_n = Wgt_4_227;
         Mult_Buf[32].Feature_n = FeatureBuf_228;
         Mult_Buf[32].Weight_n = Wgt_4_228;
         Mult_Buf[33].Feature_n = FeatureBuf_229;
         Mult_Buf[33].Weight_n = Wgt_4_229;
         Mult_Buf[34].Feature_n = FeatureBuf_230;
         Mult_Buf[34].Weight_n = Wgt_4_230;
         Mult_Buf[35].Feature_n = FeatureBuf_231;
         Mult_Buf[35].Weight_n = Wgt_4_231;
         Mult_Buf[36].Feature_n = FeatureBuf_232;
         Mult_Buf[36].Weight_n = Wgt_4_232;
         Mult_Buf[37].Feature_n = FeatureBuf_233;
         Mult_Buf[37].Weight_n = Wgt_4_233;
         Mult_Buf[38].Feature_n = FeatureBuf_234;
         Mult_Buf[38].Weight_n = Wgt_4_234;
         Mult_Buf[39].Feature_n = FeatureBuf_235;
         Mult_Buf[39].Weight_n = Wgt_4_235;
         Mult_Buf[40].Feature_n = FeatureBuf_236;
         Mult_Buf[40].Weight_n = Wgt_4_236;
         Mult_Buf[41].Feature_n = FeatureBuf_237;
         Mult_Buf[41].Weight_n = Wgt_4_237;
         Mult_Buf[42].Feature_n = FeatureBuf_238;
         Mult_Buf[42].Weight_n = Wgt_4_238;
         Mult_Buf[43].Feature_n = FeatureBuf_239;
         Mult_Buf[43].Weight_n = Wgt_4_239;
         Mult_Buf[44].Feature_n = FeatureBuf_240;
         Mult_Buf[44].Weight_n = Wgt_4_240;
         Mult_Buf[45].Feature_n = FeatureBuf_241;
         Mult_Buf[45].Weight_n = Wgt_4_241;
         Mult_Buf[46].Feature_n = FeatureBuf_242;
         Mult_Buf[46].Weight_n = Wgt_4_242;
         Mult_Buf[47].Feature_n = FeatureBuf_243;
         Mult_Buf[47].Weight_n = Wgt_4_243;
         Mult_Buf[48].Feature_n = FeatureBuf_244;
         Mult_Buf[48].Weight_n = Wgt_4_244;
         Mult_Buf[49].Feature_n = FeatureBuf_245;
         Mult_Buf[49].Weight_n = Wgt_4_245;
         Mult_Buf[50].Feature_n = FeatureBuf_246;
         Mult_Buf[50].Weight_n = Wgt_4_246;
         Mult_Buf[51].Feature_n = FeatureBuf_247;
         Mult_Buf[51].Weight_n = Wgt_4_247;
         Mult_Buf[52].Feature_n = FeatureBuf_248;
         Mult_Buf[52].Weight_n = Wgt_4_248;
         Mult_Buf[53].Feature_n = FeatureBuf_249;
         Mult_Buf[53].Weight_n = Wgt_4_249;
         Mult_Buf[54].Feature_n = FeatureBuf_250;
         Mult_Buf[54].Weight_n = Wgt_4_250;
         Mult_Buf[55].Feature_n = FeatureBuf_251;
         Mult_Buf[55].Weight_n = Wgt_4_251;
         Mult_Buf[56].Feature_n = FeatureBuf_252;
         Mult_Buf[56].Weight_n = Wgt_4_252;
         Mult_Buf[57].Feature_n = FeatureBuf_253;
         Mult_Buf[57].Weight_n = Wgt_4_253;
         Mult_Buf[58].Feature_n = FeatureBuf_254;
         Mult_Buf[58].Weight_n = Wgt_4_254;
         Mult_Buf[59].Feature_n = FeatureBuf_255;
         Mult_Buf[59].Weight_n = Wgt_4_255;
         Mult_Buf[60].Feature_n = FeatureBuf_256;
         Mult_Buf[60].Weight_n = Wgt_4_256;
         Mult_Buf[61].Feature_n = FeatureBuf_257;
         Mult_Buf[61].Weight_n = Wgt_4_257;
         Mult_Buf[62].Feature_n = FeatureBuf_258;
         Mult_Buf[62].Weight_n = Wgt_4_258;
         Mult_Buf[63].Feature_n = FeatureBuf_259;
         Mult_Buf[63].Weight_n = Wgt_4_259;
         Mult_Buf[64].Feature_n = FeatureBuf_260;
         Mult_Buf[64].Weight_n = Wgt_4_260;
         Mult_Buf[65].Feature_n = FeatureBuf_261;
         Mult_Buf[65].Weight_n = Wgt_4_261;
         Mult_Buf[66].Feature_n = FeatureBuf_262;
         Mult_Buf[66].Weight_n = Wgt_4_262;
         Mult_Buf[67].Feature_n = FeatureBuf_263;
         Mult_Buf[67].Weight_n = Wgt_4_263;
         Mult_Buf[68].Feature_n = FeatureBuf_264;
         Mult_Buf[68].Weight_n = Wgt_4_264;
         Mult_Buf[69].Feature_n = FeatureBuf_265;
         Mult_Buf[69].Weight_n = Wgt_4_265;
         Mult_Buf[70].Feature_n = FeatureBuf_266;
         Mult_Buf[70].Weight_n = Wgt_4_266;
         Mult_Buf[71].Feature_n = FeatureBuf_267;
         Mult_Buf[71].Weight_n = Wgt_4_267;
         Mult_Buf[72].Feature_n = FeatureBuf_268;
         Mult_Buf[72].Weight_n = Wgt_4_268;
         Mult_Buf[73].Feature_n = FeatureBuf_269;
         Mult_Buf[73].Weight_n = Wgt_4_269;
         Mult_Buf[74].Feature_n = FeatureBuf_270;
         Mult_Buf[74].Weight_n = Wgt_4_270;
         Mult_Buf[75].Feature_n = FeatureBuf_271;
         Mult_Buf[75].Weight_n = Wgt_4_271;
         Mult_Buf[76].Feature_n = FeatureBuf_272;
         Mult_Buf[76].Weight_n = Wgt_4_272;
         Mult_Buf[77].Feature_n = FeatureBuf_273;
         Mult_Buf[77].Weight_n = Wgt_4_273;
         Mult_Buf[78].Feature_n = FeatureBuf_274;
         Mult_Buf[78].Weight_n = Wgt_4_274;
         Mult_Buf[79].Feature_n = FeatureBuf_275;
         Mult_Buf[79].Weight_n = Wgt_4_275;
         Mult_Buf[80].Feature_n = FeatureBuf_276;
         Mult_Buf[80].Weight_n = Wgt_4_276;
         Mult_Buf[81].Feature_n = FeatureBuf_277;
         Mult_Buf[81].Weight_n = Wgt_4_277;
         Mult_Buf[82].Feature_n = FeatureBuf_278;
         Mult_Buf[82].Weight_n = Wgt_4_278;
         Mult_Buf[83].Feature_n = FeatureBuf_279;
         Mult_Buf[83].Weight_n = Wgt_4_279;
         Mult_Buf[84].Feature_n = FeatureBuf_280;
         Mult_Buf[84].Weight_n = Wgt_4_280;
         Mult_Buf[85].Feature_n = FeatureBuf_281;
         Mult_Buf[85].Weight_n = Wgt_4_281;
         Mult_Buf[86].Feature_n = FeatureBuf_282;
         Mult_Buf[86].Weight_n = Wgt_4_282;
         Mult_Buf[87].Feature_n = FeatureBuf_283;
         Mult_Buf[87].Weight_n = Wgt_4_283;
         Mult_Buf[88].Feature_n = FeatureBuf_284;
         Mult_Buf[88].Weight_n = Wgt_4_284;
         Mult_Buf[89].Feature_n = FeatureBuf_285;
         Mult_Buf[89].Weight_n = Wgt_4_285;
         Mult_Buf[90].Feature_n = FeatureBuf_286;
         Mult_Buf[90].Weight_n = Wgt_4_286;
         Mult_Buf[91].Feature_n = FeatureBuf_287;
         Mult_Buf[91].Weight_n = Wgt_4_287;
         Mult_Buf[92].Feature_n = FeatureBuf_288;
         Mult_Buf[92].Weight_n = Wgt_4_288;
         Mult_Buf[93].Feature_n = FeatureBuf_289;
         Mult_Buf[93].Weight_n = Wgt_4_289;
         Mult_Buf[94].Feature_n = FeatureBuf_290;
         Mult_Buf[94].Weight_n = Wgt_4_290;
         Mult_Buf[95].Feature_n = FeatureBuf_291;
         Mult_Buf[95].Weight_n = Wgt_4_291;
         Mult_Buf[96].Feature_n = FeatureBuf_292;
         Mult_Buf[96].Weight_n = Wgt_4_292;
         Mult_Buf[97].Feature_n = FeatureBuf_293;
         Mult_Buf[97].Weight_n = Wgt_4_293;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     //Collect Partial result form Adder
         Res_1_4_n = Part_Res;
     end
    37:begin
     nxt_state = 38;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_294;
         Mult_Buf[0].Weight_n = Wgt_4_294;
         Mult_Buf[1].Feature_n = FeatureBuf_295;
         Mult_Buf[1].Weight_n = Wgt_4_295;
         Mult_Buf[2].Feature_n = FeatureBuf_296;
         Mult_Buf[2].Weight_n = Wgt_4_296;
         Mult_Buf[3].Feature_n = FeatureBuf_297;
         Mult_Buf[3].Weight_n = Wgt_4_297;
         Mult_Buf[4].Feature_n = FeatureBuf_298;
         Mult_Buf[4].Weight_n = Wgt_4_298;
         Mult_Buf[5].Feature_n = FeatureBuf_299;
         Mult_Buf[5].Weight_n = Wgt_4_299;
         Mult_Buf[6].Feature_n = FeatureBuf_300;
         Mult_Buf[6].Weight_n = Wgt_4_300;
         Mult_Buf[7].Feature_n = FeatureBuf_301;
         Mult_Buf[7].Weight_n = Wgt_4_301;
         Mult_Buf[8].Feature_n = FeatureBuf_302;
         Mult_Buf[8].Weight_n = Wgt_4_302;
         Mult_Buf[9].Feature_n = FeatureBuf_303;
         Mult_Buf[9].Weight_n = Wgt_4_303;
         Mult_Buf[10].Feature_n = FeatureBuf_304;
         Mult_Buf[10].Weight_n = Wgt_4_304;
         Mult_Buf[11].Feature_n = FeatureBuf_305;
         Mult_Buf[11].Weight_n = Wgt_4_305;
         Mult_Buf[12].Feature_n = FeatureBuf_306;
         Mult_Buf[12].Weight_n = Wgt_4_306;
         Mult_Buf[13].Feature_n = FeatureBuf_307;
         Mult_Buf[13].Weight_n = Wgt_4_307;
         Mult_Buf[14].Feature_n = FeatureBuf_308;
         Mult_Buf[14].Weight_n = Wgt_4_308;
         Mult_Buf[15].Feature_n = FeatureBuf_309;
         Mult_Buf[15].Weight_n = Wgt_4_309;
         Mult_Buf[16].Feature_n = FeatureBuf_310;
         Mult_Buf[16].Weight_n = Wgt_4_310;
         Mult_Buf[17].Feature_n = FeatureBuf_311;
         Mult_Buf[17].Weight_n = Wgt_4_311;
         Mult_Buf[18].Feature_n = FeatureBuf_312;
         Mult_Buf[18].Weight_n = Wgt_4_312;
         Mult_Buf[19].Feature_n = FeatureBuf_313;
         Mult_Buf[19].Weight_n = Wgt_4_313;
         Mult_Buf[20].Feature_n = FeatureBuf_314;
         Mult_Buf[20].Weight_n = Wgt_4_314;
         Mult_Buf[21].Feature_n = FeatureBuf_315;
         Mult_Buf[21].Weight_n = Wgt_4_315;
         Mult_Buf[22].Feature_n = FeatureBuf_316;
         Mult_Buf[22].Weight_n = Wgt_4_316;
         Mult_Buf[23].Feature_n = FeatureBuf_317;
         Mult_Buf[23].Weight_n = Wgt_4_317;
         Mult_Buf[24].Feature_n = FeatureBuf_318;
         Mult_Buf[24].Weight_n = Wgt_4_318;
         Mult_Buf[25].Feature_n = FeatureBuf_319;
         Mult_Buf[25].Weight_n = Wgt_4_319;
         Mult_Buf[26].Feature_n = FeatureBuf_320;
         Mult_Buf[26].Weight_n = Wgt_4_320;
         Mult_Buf[27].Feature_n = FeatureBuf_321;
         Mult_Buf[27].Weight_n = Wgt_4_321;
         Mult_Buf[28].Feature_n = FeatureBuf_322;
         Mult_Buf[28].Weight_n = Wgt_4_322;
         Mult_Buf[29].Feature_n = FeatureBuf_323;
         Mult_Buf[29].Weight_n = Wgt_4_323;
         Mult_Buf[30].Feature_n = FeatureBuf_324;
         Mult_Buf[30].Weight_n = Wgt_4_324;
         Mult_Buf[31].Feature_n = FeatureBuf_325;
         Mult_Buf[31].Weight_n = Wgt_4_325;
         Mult_Buf[32].Feature_n = FeatureBuf_326;
         Mult_Buf[32].Weight_n = Wgt_4_326;
         Mult_Buf[33].Feature_n = FeatureBuf_327;
         Mult_Buf[33].Weight_n = Wgt_4_327;
         Mult_Buf[34].Feature_n = FeatureBuf_328;
         Mult_Buf[34].Weight_n = Wgt_4_328;
         Mult_Buf[35].Feature_n = FeatureBuf_329;
         Mult_Buf[35].Weight_n = Wgt_4_329;
         Mult_Buf[36].Feature_n = FeatureBuf_330;
         Mult_Buf[36].Weight_n = Wgt_4_330;
         Mult_Buf[37].Feature_n = FeatureBuf_331;
         Mult_Buf[37].Weight_n = Wgt_4_331;
         Mult_Buf[38].Feature_n = FeatureBuf_332;
         Mult_Buf[38].Weight_n = Wgt_4_332;
         Mult_Buf[39].Feature_n = FeatureBuf_333;
         Mult_Buf[39].Weight_n = Wgt_4_333;
         Mult_Buf[40].Feature_n = FeatureBuf_334;
         Mult_Buf[40].Weight_n = Wgt_4_334;
         Mult_Buf[41].Feature_n = FeatureBuf_335;
         Mult_Buf[41].Weight_n = Wgt_4_335;
         Mult_Buf[42].Feature_n = FeatureBuf_336;
         Mult_Buf[42].Weight_n = Wgt_4_336;
         Mult_Buf[43].Feature_n = FeatureBuf_337;
         Mult_Buf[43].Weight_n = Wgt_4_337;
         Mult_Buf[44].Feature_n = FeatureBuf_338;
         Mult_Buf[44].Weight_n = Wgt_4_338;
         Mult_Buf[45].Feature_n = FeatureBuf_339;
         Mult_Buf[45].Weight_n = Wgt_4_339;
         Mult_Buf[46].Feature_n = FeatureBuf_340;
         Mult_Buf[46].Weight_n = Wgt_4_340;
         Mult_Buf[47].Feature_n = FeatureBuf_341;
         Mult_Buf[47].Weight_n = Wgt_4_341;
         Mult_Buf[48].Feature_n = FeatureBuf_342;
         Mult_Buf[48].Weight_n = Wgt_4_342;
         Mult_Buf[49].Feature_n = FeatureBuf_343;
         Mult_Buf[49].Weight_n = Wgt_4_343;
         Mult_Buf[50].Feature_n = FeatureBuf_344;
         Mult_Buf[50].Weight_n = Wgt_4_344;
         Mult_Buf[51].Feature_n = FeatureBuf_345;
         Mult_Buf[51].Weight_n = Wgt_4_345;
         Mult_Buf[52].Feature_n = FeatureBuf_346;
         Mult_Buf[52].Weight_n = Wgt_4_346;
         Mult_Buf[53].Feature_n = FeatureBuf_347;
         Mult_Buf[53].Weight_n = Wgt_4_347;
         Mult_Buf[54].Feature_n = FeatureBuf_348;
         Mult_Buf[54].Weight_n = Wgt_4_348;
         Mult_Buf[55].Feature_n = FeatureBuf_349;
         Mult_Buf[55].Weight_n = Wgt_4_349;
         Mult_Buf[56].Feature_n = FeatureBuf_350;
         Mult_Buf[56].Weight_n = Wgt_4_350;
         Mult_Buf[57].Feature_n = FeatureBuf_351;
         Mult_Buf[57].Weight_n = Wgt_4_351;
         Mult_Buf[58].Feature_n = FeatureBuf_352;
         Mult_Buf[58].Weight_n = Wgt_4_352;
         Mult_Buf[59].Feature_n = FeatureBuf_353;
         Mult_Buf[59].Weight_n = Wgt_4_353;
         Mult_Buf[60].Feature_n = FeatureBuf_354;
         Mult_Buf[60].Weight_n = Wgt_4_354;
         Mult_Buf[61].Feature_n = FeatureBuf_355;
         Mult_Buf[61].Weight_n = Wgt_4_355;
         Mult_Buf[62].Feature_n = FeatureBuf_356;
         Mult_Buf[62].Weight_n = Wgt_4_356;
         Mult_Buf[63].Feature_n = FeatureBuf_357;
         Mult_Buf[63].Weight_n = Wgt_4_357;
         Mult_Buf[64].Feature_n = FeatureBuf_358;
         Mult_Buf[64].Weight_n = Wgt_4_358;
         Mult_Buf[65].Feature_n = FeatureBuf_359;
         Mult_Buf[65].Weight_n = Wgt_4_359;
         Mult_Buf[66].Feature_n = FeatureBuf_360;
         Mult_Buf[66].Weight_n = Wgt_4_360;
         Mult_Buf[67].Feature_n = FeatureBuf_361;
         Mult_Buf[67].Weight_n = Wgt_4_361;
         Mult_Buf[68].Feature_n = FeatureBuf_362;
         Mult_Buf[68].Weight_n = Wgt_4_362;
         Mult_Buf[69].Feature_n = FeatureBuf_363;
         Mult_Buf[69].Weight_n = Wgt_4_363;
         Mult_Buf[70].Feature_n = FeatureBuf_364;
         Mult_Buf[70].Weight_n = Wgt_4_364;
         Mult_Buf[71].Feature_n = FeatureBuf_365;
         Mult_Buf[71].Weight_n = Wgt_4_365;
         Mult_Buf[72].Feature_n = FeatureBuf_366;
         Mult_Buf[72].Weight_n = Wgt_4_366;
         Mult_Buf[73].Feature_n = FeatureBuf_367;
         Mult_Buf[73].Weight_n = Wgt_4_367;
         Mult_Buf[74].Feature_n = FeatureBuf_368;
         Mult_Buf[74].Weight_n = Wgt_4_368;
         Mult_Buf[75].Feature_n = FeatureBuf_369;
         Mult_Buf[75].Weight_n = Wgt_4_369;
         Mult_Buf[76].Feature_n = FeatureBuf_370;
         Mult_Buf[76].Weight_n = Wgt_4_370;
         Mult_Buf[77].Feature_n = FeatureBuf_371;
         Mult_Buf[77].Weight_n = Wgt_4_371;
         Mult_Buf[78].Feature_n = FeatureBuf_372;
         Mult_Buf[78].Weight_n = Wgt_4_372;
         Mult_Buf[79].Feature_n = FeatureBuf_373;
         Mult_Buf[79].Weight_n = Wgt_4_373;
         Mult_Buf[80].Feature_n = FeatureBuf_374;
         Mult_Buf[80].Weight_n = Wgt_4_374;
         Mult_Buf[81].Feature_n = FeatureBuf_375;
         Mult_Buf[81].Weight_n = Wgt_4_375;
         Mult_Buf[82].Feature_n = FeatureBuf_376;
         Mult_Buf[82].Weight_n = Wgt_4_376;
         Mult_Buf[83].Feature_n = FeatureBuf_377;
         Mult_Buf[83].Weight_n = Wgt_4_377;
         Mult_Buf[84].Feature_n = FeatureBuf_378;
         Mult_Buf[84].Weight_n = Wgt_4_378;
         Mult_Buf[85].Feature_n = FeatureBuf_379;
         Mult_Buf[85].Weight_n = Wgt_4_379;
         Mult_Buf[86].Feature_n = FeatureBuf_380;
         Mult_Buf[86].Weight_n = Wgt_4_380;
         Mult_Buf[87].Feature_n = FeatureBuf_381;
         Mult_Buf[87].Weight_n = Wgt_4_381;
         Mult_Buf[88].Feature_n = FeatureBuf_382;
         Mult_Buf[88].Weight_n = Wgt_4_382;
         Mult_Buf[89].Feature_n = FeatureBuf_383;
         Mult_Buf[89].Weight_n = Wgt_4_383;
         Mult_Buf[90].Feature_n = FeatureBuf_384;
         Mult_Buf[90].Weight_n = Wgt_4_384;
         Mult_Buf[91].Feature_n = FeatureBuf_385;
         Mult_Buf[91].Weight_n = Wgt_4_385;
         Mult_Buf[92].Feature_n = FeatureBuf_386;
         Mult_Buf[92].Weight_n = Wgt_4_386;
         Mult_Buf[93].Feature_n = FeatureBuf_387;
         Mult_Buf[93].Weight_n = Wgt_4_387;
         Mult_Buf[94].Feature_n = FeatureBuf_388;
         Mult_Buf[94].Weight_n = Wgt_4_388;
         Mult_Buf[95].Feature_n = FeatureBuf_389;
         Mult_Buf[95].Weight_n = Wgt_4_389;
         Mult_Buf[96].Feature_n = FeatureBuf_390;
         Mult_Buf[96].Weight_n = Wgt_4_390;
         Mult_Buf[97].Feature_n = FeatureBuf_391;
         Mult_Buf[97].Weight_n = Wgt_4_391;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     //Collect Partial result form Adder
         Res_1_5_n = Part_Res;
     //Collect result from final Adder
         Res0_n = Final_Res;
     end
    38:begin
     nxt_state = 39;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_392;
         Mult_Buf[0].Weight_n = Wgt_4_392;
         Mult_Buf[1].Feature_n = FeatureBuf_393;
         Mult_Buf[1].Weight_n = Wgt_4_393;
         Mult_Buf[2].Feature_n = FeatureBuf_394;
         Mult_Buf[2].Weight_n = Wgt_4_394;
         Mult_Buf[3].Feature_n = FeatureBuf_395;
         Mult_Buf[3].Weight_n = Wgt_4_395;
         Mult_Buf[4].Feature_n = FeatureBuf_396;
         Mult_Buf[4].Weight_n = Wgt_4_396;
         Mult_Buf[5].Feature_n = FeatureBuf_397;
         Mult_Buf[5].Weight_n = Wgt_4_397;
         Mult_Buf[6].Feature_n = FeatureBuf_398;
         Mult_Buf[6].Weight_n = Wgt_4_398;
         Mult_Buf[7].Feature_n = FeatureBuf_399;
         Mult_Buf[7].Weight_n = Wgt_4_399;
         Mult_Buf[8].Feature_n = FeatureBuf_400;
         Mult_Buf[8].Weight_n = Wgt_4_400;
         Mult_Buf[9].Feature_n = FeatureBuf_401;
         Mult_Buf[9].Weight_n = Wgt_4_401;
         Mult_Buf[10].Feature_n = FeatureBuf_402;
         Mult_Buf[10].Weight_n = Wgt_4_402;
         Mult_Buf[11].Feature_n = FeatureBuf_403;
         Mult_Buf[11].Weight_n = Wgt_4_403;
         Mult_Buf[12].Feature_n = FeatureBuf_404;
         Mult_Buf[12].Weight_n = Wgt_4_404;
         Mult_Buf[13].Feature_n = FeatureBuf_405;
         Mult_Buf[13].Weight_n = Wgt_4_405;
         Mult_Buf[14].Feature_n = FeatureBuf_406;
         Mult_Buf[14].Weight_n = Wgt_4_406;
         Mult_Buf[15].Feature_n = FeatureBuf_407;
         Mult_Buf[15].Weight_n = Wgt_4_407;
         Mult_Buf[16].Feature_n = FeatureBuf_408;
         Mult_Buf[16].Weight_n = Wgt_4_408;
         Mult_Buf[17].Feature_n = FeatureBuf_409;
         Mult_Buf[17].Weight_n = Wgt_4_409;
         Mult_Buf[18].Feature_n = FeatureBuf_410;
         Mult_Buf[18].Weight_n = Wgt_4_410;
         Mult_Buf[19].Feature_n = FeatureBuf_411;
         Mult_Buf[19].Weight_n = Wgt_4_411;
         Mult_Buf[20].Feature_n = FeatureBuf_412;
         Mult_Buf[20].Weight_n = Wgt_4_412;
         Mult_Buf[21].Feature_n = FeatureBuf_413;
         Mult_Buf[21].Weight_n = Wgt_4_413;
         Mult_Buf[22].Feature_n = FeatureBuf_414;
         Mult_Buf[22].Weight_n = Wgt_4_414;
         Mult_Buf[23].Feature_n = FeatureBuf_415;
         Mult_Buf[23].Weight_n = Wgt_4_415;
         Mult_Buf[24].Feature_n = FeatureBuf_416;
         Mult_Buf[24].Weight_n = Wgt_4_416;
         Mult_Buf[25].Feature_n = FeatureBuf_417;
         Mult_Buf[25].Weight_n = Wgt_4_417;
         Mult_Buf[26].Feature_n = FeatureBuf_418;
         Mult_Buf[26].Weight_n = Wgt_4_418;
         Mult_Buf[27].Feature_n = FeatureBuf_419;
         Mult_Buf[27].Weight_n = Wgt_4_419;
         Mult_Buf[28].Feature_n = FeatureBuf_420;
         Mult_Buf[28].Weight_n = Wgt_4_420;
         Mult_Buf[29].Feature_n = FeatureBuf_421;
         Mult_Buf[29].Weight_n = Wgt_4_421;
         Mult_Buf[30].Feature_n = FeatureBuf_422;
         Mult_Buf[30].Weight_n = Wgt_4_422;
         Mult_Buf[31].Feature_n = FeatureBuf_423;
         Mult_Buf[31].Weight_n = Wgt_4_423;
         Mult_Buf[32].Feature_n = FeatureBuf_424;
         Mult_Buf[32].Weight_n = Wgt_4_424;
         Mult_Buf[33].Feature_n = FeatureBuf_425;
         Mult_Buf[33].Weight_n = Wgt_4_425;
         Mult_Buf[34].Feature_n = FeatureBuf_426;
         Mult_Buf[34].Weight_n = Wgt_4_426;
         Mult_Buf[35].Feature_n = FeatureBuf_427;
         Mult_Buf[35].Weight_n = Wgt_4_427;
         Mult_Buf[36].Feature_n = FeatureBuf_428;
         Mult_Buf[36].Weight_n = Wgt_4_428;
         Mult_Buf[37].Feature_n = FeatureBuf_429;
         Mult_Buf[37].Weight_n = Wgt_4_429;
         Mult_Buf[38].Feature_n = FeatureBuf_430;
         Mult_Buf[38].Weight_n = Wgt_4_430;
         Mult_Buf[39].Feature_n = FeatureBuf_431;
         Mult_Buf[39].Weight_n = Wgt_4_431;
         Mult_Buf[40].Feature_n = FeatureBuf_432;
         Mult_Buf[40].Weight_n = Wgt_4_432;
         Mult_Buf[41].Feature_n = FeatureBuf_433;
         Mult_Buf[41].Weight_n = Wgt_4_433;
         Mult_Buf[42].Feature_n = FeatureBuf_434;
         Mult_Buf[42].Weight_n = Wgt_4_434;
         Mult_Buf[43].Feature_n = FeatureBuf_435;
         Mult_Buf[43].Weight_n = Wgt_4_435;
         Mult_Buf[44].Feature_n = FeatureBuf_436;
         Mult_Buf[44].Weight_n = Wgt_4_436;
         Mult_Buf[45].Feature_n = FeatureBuf_437;
         Mult_Buf[45].Weight_n = Wgt_4_437;
         Mult_Buf[46].Feature_n = FeatureBuf_438;
         Mult_Buf[46].Weight_n = Wgt_4_438;
         Mult_Buf[47].Feature_n = FeatureBuf_439;
         Mult_Buf[47].Weight_n = Wgt_4_439;
         Mult_Buf[48].Feature_n = FeatureBuf_440;
         Mult_Buf[48].Weight_n = Wgt_4_440;
         Mult_Buf[49].Feature_n = FeatureBuf_441;
         Mult_Buf[49].Weight_n = Wgt_4_441;
         Mult_Buf[50].Feature_n = FeatureBuf_442;
         Mult_Buf[50].Weight_n = Wgt_4_442;
         Mult_Buf[51].Feature_n = FeatureBuf_443;
         Mult_Buf[51].Weight_n = Wgt_4_443;
         Mult_Buf[52].Feature_n = FeatureBuf_444;
         Mult_Buf[52].Weight_n = Wgt_4_444;
         Mult_Buf[53].Feature_n = FeatureBuf_445;
         Mult_Buf[53].Weight_n = Wgt_4_445;
         Mult_Buf[54].Feature_n = FeatureBuf_446;
         Mult_Buf[54].Weight_n = Wgt_4_446;
         Mult_Buf[55].Feature_n = FeatureBuf_447;
         Mult_Buf[55].Weight_n = Wgt_4_447;
         Mult_Buf[56].Feature_n = FeatureBuf_448;
         Mult_Buf[56].Weight_n = Wgt_4_448;
         Mult_Buf[57].Feature_n = FeatureBuf_449;
         Mult_Buf[57].Weight_n = Wgt_4_449;
         Mult_Buf[58].Feature_n = FeatureBuf_450;
         Mult_Buf[58].Weight_n = Wgt_4_450;
         Mult_Buf[59].Feature_n = FeatureBuf_451;
         Mult_Buf[59].Weight_n = Wgt_4_451;
         Mult_Buf[60].Feature_n = FeatureBuf_452;
         Mult_Buf[60].Weight_n = Wgt_4_452;
         Mult_Buf[61].Feature_n = FeatureBuf_453;
         Mult_Buf[61].Weight_n = Wgt_4_453;
         Mult_Buf[62].Feature_n = FeatureBuf_454;
         Mult_Buf[62].Weight_n = Wgt_4_454;
         Mult_Buf[63].Feature_n = FeatureBuf_455;
         Mult_Buf[63].Weight_n = Wgt_4_455;
         Mult_Buf[64].Feature_n = FeatureBuf_456;
         Mult_Buf[64].Weight_n = Wgt_4_456;
         Mult_Buf[65].Feature_n = FeatureBuf_457;
         Mult_Buf[65].Weight_n = Wgt_4_457;
         Mult_Buf[66].Feature_n = FeatureBuf_458;
         Mult_Buf[66].Weight_n = Wgt_4_458;
         Mult_Buf[67].Feature_n = FeatureBuf_459;
         Mult_Buf[67].Weight_n = Wgt_4_459;
         Mult_Buf[68].Feature_n = FeatureBuf_460;
         Mult_Buf[68].Weight_n = Wgt_4_460;
         Mult_Buf[69].Feature_n = FeatureBuf_461;
         Mult_Buf[69].Weight_n = Wgt_4_461;
         Mult_Buf[70].Feature_n = FeatureBuf_462;
         Mult_Buf[70].Weight_n = Wgt_4_462;
         Mult_Buf[71].Feature_n = FeatureBuf_463;
         Mult_Buf[71].Weight_n = Wgt_4_463;
         Mult_Buf[72].Feature_n = FeatureBuf_464;
         Mult_Buf[72].Weight_n = Wgt_4_464;
         Mult_Buf[73].Feature_n = FeatureBuf_465;
         Mult_Buf[73].Weight_n = Wgt_4_465;
         Mult_Buf[74].Feature_n = FeatureBuf_466;
         Mult_Buf[74].Weight_n = Wgt_4_466;
         Mult_Buf[75].Feature_n = FeatureBuf_467;
         Mult_Buf[75].Weight_n = Wgt_4_467;
         Mult_Buf[76].Feature_n = FeatureBuf_468;
         Mult_Buf[76].Weight_n = Wgt_4_468;
         Mult_Buf[77].Feature_n = FeatureBuf_469;
         Mult_Buf[77].Weight_n = Wgt_4_469;
         Mult_Buf[78].Feature_n = FeatureBuf_470;
         Mult_Buf[78].Weight_n = Wgt_4_470;
         Mult_Buf[79].Feature_n = FeatureBuf_471;
         Mult_Buf[79].Weight_n = Wgt_4_471;
         Mult_Buf[80].Feature_n = FeatureBuf_472;
         Mult_Buf[80].Weight_n = Wgt_4_472;
         Mult_Buf[81].Feature_n = FeatureBuf_473;
         Mult_Buf[81].Weight_n = Wgt_4_473;
         Mult_Buf[82].Feature_n = FeatureBuf_474;
         Mult_Buf[82].Weight_n = Wgt_4_474;
         Mult_Buf[83].Feature_n = FeatureBuf_475;
         Mult_Buf[83].Weight_n = Wgt_4_475;
         Mult_Buf[84].Feature_n = FeatureBuf_476;
         Mult_Buf[84].Weight_n = Wgt_4_476;
         Mult_Buf[85].Feature_n = FeatureBuf_477;
         Mult_Buf[85].Weight_n = Wgt_4_477;
         Mult_Buf[86].Feature_n = FeatureBuf_478;
         Mult_Buf[86].Weight_n = Wgt_4_478;
         Mult_Buf[87].Feature_n = FeatureBuf_479;
         Mult_Buf[87].Weight_n = Wgt_4_479;
         Mult_Buf[88].Feature_n = FeatureBuf_480;
         Mult_Buf[88].Weight_n = Wgt_4_480;
         Mult_Buf[89].Feature_n = FeatureBuf_481;
         Mult_Buf[89].Weight_n = Wgt_4_481;
         Mult_Buf[90].Feature_n = FeatureBuf_482;
         Mult_Buf[90].Weight_n = Wgt_4_482;
         Mult_Buf[91].Feature_n = FeatureBuf_483;
         Mult_Buf[91].Weight_n = Wgt_4_483;
         Mult_Buf[92].Feature_n = FeatureBuf_484;
         Mult_Buf[92].Weight_n = Wgt_4_484;
         Mult_Buf[93].Feature_n = FeatureBuf_485;
         Mult_Buf[93].Weight_n = Wgt_4_485;
         Mult_Buf[94].Feature_n = FeatureBuf_486;
         Mult_Buf[94].Weight_n = Wgt_4_486;
         Mult_Buf[95].Feature_n = FeatureBuf_487;
         Mult_Buf[95].Weight_n = Wgt_4_487;
         Mult_Buf[96].Feature_n = FeatureBuf_488;
         Mult_Buf[96].Weight_n = Wgt_4_488;
         Mult_Buf[97].Feature_n = FeatureBuf_489;
         Mult_Buf[97].Weight_n = Wgt_4_489;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     //Collect Partial result form Adder
         Res_1_6_n = Part_Res;
     end
    39:begin
     nxt_state = 40;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_490;
         Mult_Buf[0].Weight_n = Wgt_4_490;
         Mult_Buf[1].Feature_n = FeatureBuf_491;
         Mult_Buf[1].Weight_n = Wgt_4_491;
         Mult_Buf[2].Feature_n = FeatureBuf_492;
         Mult_Buf[2].Weight_n = Wgt_4_492;
         Mult_Buf[3].Feature_n = FeatureBuf_493;
         Mult_Buf[3].Weight_n = Wgt_4_493;
         Mult_Buf[4].Feature_n = FeatureBuf_494;
         Mult_Buf[4].Weight_n = Wgt_4_494;
         Mult_Buf[5].Feature_n = FeatureBuf_495;
         Mult_Buf[5].Weight_n = Wgt_4_495;
         Mult_Buf[6].Feature_n = FeatureBuf_496;
         Mult_Buf[6].Weight_n = Wgt_4_496;
         Mult_Buf[7].Feature_n = FeatureBuf_497;
         Mult_Buf[7].Weight_n = Wgt_4_497;
         Mult_Buf[8].Feature_n = FeatureBuf_498;
         Mult_Buf[8].Weight_n = Wgt_4_498;
         Mult_Buf[9].Feature_n = FeatureBuf_499;
         Mult_Buf[9].Weight_n = Wgt_4_499;
         Mult_Buf[10].Feature_n = FeatureBuf_500;
         Mult_Buf[10].Weight_n = Wgt_4_500;
         Mult_Buf[11].Feature_n = FeatureBuf_501;
         Mult_Buf[11].Weight_n = Wgt_4_501;
         Mult_Buf[12].Feature_n = FeatureBuf_502;
         Mult_Buf[12].Weight_n = Wgt_4_502;
         Mult_Buf[13].Feature_n = FeatureBuf_503;
         Mult_Buf[13].Weight_n = Wgt_4_503;
         Mult_Buf[14].Feature_n = FeatureBuf_504;
         Mult_Buf[14].Weight_n = Wgt_4_504;
         Mult_Buf[15].Feature_n = FeatureBuf_505;
         Mult_Buf[15].Weight_n = Wgt_4_505;
         Mult_Buf[16].Feature_n = FeatureBuf_506;
         Mult_Buf[16].Weight_n = Wgt_4_506;
         Mult_Buf[17].Feature_n = FeatureBuf_507;
         Mult_Buf[17].Weight_n = Wgt_4_507;
         Mult_Buf[18].Feature_n = FeatureBuf_508;
         Mult_Buf[18].Weight_n = Wgt_4_508;
         Mult_Buf[19].Feature_n = FeatureBuf_509;
         Mult_Buf[19].Weight_n = Wgt_4_509;
         Mult_Buf[20].Feature_n = FeatureBuf_510;
         Mult_Buf[20].Weight_n = Wgt_4_510;
         Mult_Buf[21].Feature_n = FeatureBuf_511;
         Mult_Buf[21].Weight_n = Wgt_4_511;
         Mult_Buf[22].Feature_n = FeatureBuf_512;
         Mult_Buf[22].Weight_n = Wgt_4_512;
         Mult_Buf[23].Feature_n = FeatureBuf_513;
         Mult_Buf[23].Weight_n = Wgt_4_513;
         Mult_Buf[24].Feature_n = FeatureBuf_514;
         Mult_Buf[24].Weight_n = Wgt_4_514;
         Mult_Buf[25].Feature_n = FeatureBuf_515;
         Mult_Buf[25].Weight_n = Wgt_4_515;
         Mult_Buf[26].Feature_n = FeatureBuf_516;
         Mult_Buf[26].Weight_n = Wgt_4_516;
         Mult_Buf[27].Feature_n = FeatureBuf_517;
         Mult_Buf[27].Weight_n = Wgt_4_517;
         Mult_Buf[28].Feature_n = FeatureBuf_518;
         Mult_Buf[28].Weight_n = Wgt_4_518;
         Mult_Buf[29].Feature_n = FeatureBuf_519;
         Mult_Buf[29].Weight_n = Wgt_4_519;
         Mult_Buf[30].Feature_n = FeatureBuf_520;
         Mult_Buf[30].Weight_n = Wgt_4_520;
         Mult_Buf[31].Feature_n = FeatureBuf_521;
         Mult_Buf[31].Weight_n = Wgt_4_521;
         Mult_Buf[32].Feature_n = FeatureBuf_522;
         Mult_Buf[32].Weight_n = Wgt_4_522;
         Mult_Buf[33].Feature_n = FeatureBuf_523;
         Mult_Buf[33].Weight_n = Wgt_4_523;
         Mult_Buf[34].Feature_n = FeatureBuf_524;
         Mult_Buf[34].Weight_n = Wgt_4_524;
         Mult_Buf[35].Feature_n = FeatureBuf_525;
         Mult_Buf[35].Weight_n = Wgt_4_525;
         Mult_Buf[36].Feature_n = FeatureBuf_526;
         Mult_Buf[36].Weight_n = Wgt_4_526;
         Mult_Buf[37].Feature_n = FeatureBuf_527;
         Mult_Buf[37].Weight_n = Wgt_4_527;
         Mult_Buf[38].Feature_n = FeatureBuf_528;
         Mult_Buf[38].Weight_n = Wgt_4_528;
         Mult_Buf[39].Feature_n = FeatureBuf_529;
         Mult_Buf[39].Weight_n = Wgt_4_529;
         Mult_Buf[40].Feature_n = FeatureBuf_530;
         Mult_Buf[40].Weight_n = Wgt_4_530;
         Mult_Buf[41].Feature_n = FeatureBuf_531;
         Mult_Buf[41].Weight_n = Wgt_4_531;
         Mult_Buf[42].Feature_n = FeatureBuf_532;
         Mult_Buf[42].Weight_n = Wgt_4_532;
         Mult_Buf[43].Feature_n = FeatureBuf_533;
         Mult_Buf[43].Weight_n = Wgt_4_533;
         Mult_Buf[44].Feature_n = FeatureBuf_534;
         Mult_Buf[44].Weight_n = Wgt_4_534;
         Mult_Buf[45].Feature_n = FeatureBuf_535;
         Mult_Buf[45].Weight_n = Wgt_4_535;
         Mult_Buf[46].Feature_n = FeatureBuf_536;
         Mult_Buf[46].Weight_n = Wgt_4_536;
         Mult_Buf[47].Feature_n = FeatureBuf_537;
         Mult_Buf[47].Weight_n = Wgt_4_537;
         Mult_Buf[48].Feature_n = FeatureBuf_538;
         Mult_Buf[48].Weight_n = Wgt_4_538;
         Mult_Buf[49].Feature_n = FeatureBuf_539;
         Mult_Buf[49].Weight_n = Wgt_4_539;
         Mult_Buf[50].Feature_n = FeatureBuf_540;
         Mult_Buf[50].Weight_n = Wgt_4_540;
         Mult_Buf[51].Feature_n = FeatureBuf_541;
         Mult_Buf[51].Weight_n = Wgt_4_541;
         Mult_Buf[52].Feature_n = FeatureBuf_542;
         Mult_Buf[52].Weight_n = Wgt_4_542;
         Mult_Buf[53].Feature_n = FeatureBuf_543;
         Mult_Buf[53].Weight_n = Wgt_4_543;
         Mult_Buf[54].Feature_n = FeatureBuf_544;
         Mult_Buf[54].Weight_n = Wgt_4_544;
         Mult_Buf[55].Feature_n = FeatureBuf_545;
         Mult_Buf[55].Weight_n = Wgt_4_545;
         Mult_Buf[56].Feature_n = FeatureBuf_546;
         Mult_Buf[56].Weight_n = Wgt_4_546;
         Mult_Buf[57].Feature_n = FeatureBuf_547;
         Mult_Buf[57].Weight_n = Wgt_4_547;
         Mult_Buf[58].Feature_n = FeatureBuf_548;
         Mult_Buf[58].Weight_n = Wgt_4_548;
         Mult_Buf[59].Feature_n = FeatureBuf_549;
         Mult_Buf[59].Weight_n = Wgt_4_549;
         Mult_Buf[60].Feature_n = FeatureBuf_550;
         Mult_Buf[60].Weight_n = Wgt_4_550;
         Mult_Buf[61].Feature_n = FeatureBuf_551;
         Mult_Buf[61].Weight_n = Wgt_4_551;
         Mult_Buf[62].Feature_n = FeatureBuf_552;
         Mult_Buf[62].Weight_n = Wgt_4_552;
         Mult_Buf[63].Feature_n = FeatureBuf_553;
         Mult_Buf[63].Weight_n = Wgt_4_553;
         Mult_Buf[64].Feature_n = FeatureBuf_554;
         Mult_Buf[64].Weight_n = Wgt_4_554;
         Mult_Buf[65].Feature_n = FeatureBuf_555;
         Mult_Buf[65].Weight_n = Wgt_4_555;
         Mult_Buf[66].Feature_n = FeatureBuf_556;
         Mult_Buf[66].Weight_n = Wgt_4_556;
         Mult_Buf[67].Feature_n = FeatureBuf_557;
         Mult_Buf[67].Weight_n = Wgt_4_557;
         Mult_Buf[68].Feature_n = FeatureBuf_558;
         Mult_Buf[68].Weight_n = Wgt_4_558;
         Mult_Buf[69].Feature_n = FeatureBuf_559;
         Mult_Buf[69].Weight_n = Wgt_4_559;
         Mult_Buf[70].Feature_n = FeatureBuf_560;
         Mult_Buf[70].Weight_n = Wgt_4_560;
         Mult_Buf[71].Feature_n = FeatureBuf_561;
         Mult_Buf[71].Weight_n = Wgt_4_561;
         Mult_Buf[72].Feature_n = FeatureBuf_562;
         Mult_Buf[72].Weight_n = Wgt_4_562;
         Mult_Buf[73].Feature_n = FeatureBuf_563;
         Mult_Buf[73].Weight_n = Wgt_4_563;
         Mult_Buf[74].Feature_n = FeatureBuf_564;
         Mult_Buf[74].Weight_n = Wgt_4_564;
         Mult_Buf[75].Feature_n = FeatureBuf_565;
         Mult_Buf[75].Weight_n = Wgt_4_565;
         Mult_Buf[76].Feature_n = FeatureBuf_566;
         Mult_Buf[76].Weight_n = Wgt_4_566;
         Mult_Buf[77].Feature_n = FeatureBuf_567;
         Mult_Buf[77].Weight_n = Wgt_4_567;
         Mult_Buf[78].Feature_n = FeatureBuf_568;
         Mult_Buf[78].Weight_n = Wgt_4_568;
         Mult_Buf[79].Feature_n = FeatureBuf_569;
         Mult_Buf[79].Weight_n = Wgt_4_569;
         Mult_Buf[80].Feature_n = FeatureBuf_570;
         Mult_Buf[80].Weight_n = Wgt_4_570;
         Mult_Buf[81].Feature_n = FeatureBuf_571;
         Mult_Buf[81].Weight_n = Wgt_4_571;
         Mult_Buf[82].Feature_n = FeatureBuf_572;
         Mult_Buf[82].Weight_n = Wgt_4_572;
         Mult_Buf[83].Feature_n = FeatureBuf_573;
         Mult_Buf[83].Weight_n = Wgt_4_573;
         Mult_Buf[84].Feature_n = FeatureBuf_574;
         Mult_Buf[84].Weight_n = Wgt_4_574;
         Mult_Buf[85].Feature_n = FeatureBuf_575;
         Mult_Buf[85].Weight_n = Wgt_4_575;
         Mult_Buf[86].Feature_n = FeatureBuf_576;
         Mult_Buf[86].Weight_n = Wgt_4_576;
         Mult_Buf[87].Feature_n = FeatureBuf_577;
         Mult_Buf[87].Weight_n = Wgt_4_577;
         Mult_Buf[88].Feature_n = FeatureBuf_578;
         Mult_Buf[88].Weight_n = Wgt_4_578;
         Mult_Buf[89].Feature_n = FeatureBuf_579;
         Mult_Buf[89].Weight_n = Wgt_4_579;
         Mult_Buf[90].Feature_n = FeatureBuf_580;
         Mult_Buf[90].Weight_n = Wgt_4_580;
         Mult_Buf[91].Feature_n = FeatureBuf_581;
         Mult_Buf[91].Weight_n = Wgt_4_581;
         Mult_Buf[92].Feature_n = FeatureBuf_582;
         Mult_Buf[92].Weight_n = Wgt_4_582;
         Mult_Buf[93].Feature_n = FeatureBuf_583;
         Mult_Buf[93].Weight_n = Wgt_4_583;
         Mult_Buf[94].Feature_n = FeatureBuf_584;
         Mult_Buf[94].Weight_n = Wgt_4_584;
         Mult_Buf[95].Feature_n = FeatureBuf_585;
         Mult_Buf[95].Weight_n = Wgt_4_585;
         Mult_Buf[96].Feature_n = FeatureBuf_586;
         Mult_Buf[96].Weight_n = Wgt_4_586;
         Mult_Buf[97].Feature_n = FeatureBuf_587;
         Mult_Buf[97].Weight_n = Wgt_4_587;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     //Collect Partial result form Adder
         Res_1_7_n = Part_Res;
     //Feed to final Adder
         A1 = Part_Res;
         A2 = Res_1_6_n;
         A3 = Res_1_5_n;
         A4 = Res_1_4_n;
         A5 = Res_1_3_n;
         A6 = Res_1_2_n;
         A7 = Res_1_1_n;
         A8 = Res_1_0_n;
     end
    40:begin
     nxt_state = 41;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_588;
         Mult_Buf[0].Weight_n = Wgt_4_588;
         Mult_Buf[1].Feature_n = FeatureBuf_589;
         Mult_Buf[1].Weight_n = Wgt_4_589;
         Mult_Buf[2].Feature_n = FeatureBuf_590;
         Mult_Buf[2].Weight_n = Wgt_4_590;
         Mult_Buf[3].Feature_n = FeatureBuf_591;
         Mult_Buf[3].Weight_n = Wgt_4_591;
         Mult_Buf[4].Feature_n = FeatureBuf_592;
         Mult_Buf[4].Weight_n = Wgt_4_592;
         Mult_Buf[5].Feature_n = FeatureBuf_593;
         Mult_Buf[5].Weight_n = Wgt_4_593;
         Mult_Buf[6].Feature_n = FeatureBuf_594;
         Mult_Buf[6].Weight_n = Wgt_4_594;
         Mult_Buf[7].Feature_n = FeatureBuf_595;
         Mult_Buf[7].Weight_n = Wgt_4_595;
         Mult_Buf[8].Feature_n = FeatureBuf_596;
         Mult_Buf[8].Weight_n = Wgt_4_596;
         Mult_Buf[9].Feature_n = FeatureBuf_597;
         Mult_Buf[9].Weight_n = Wgt_4_597;
         Mult_Buf[10].Feature_n = FeatureBuf_598;
         Mult_Buf[10].Weight_n = Wgt_4_598;
         Mult_Buf[11].Feature_n = FeatureBuf_599;
         Mult_Buf[11].Weight_n = Wgt_4_599;
         Mult_Buf[12].Feature_n = FeatureBuf_600;
         Mult_Buf[12].Weight_n = Wgt_4_600;
         Mult_Buf[13].Feature_n = FeatureBuf_601;
         Mult_Buf[13].Weight_n = Wgt_4_601;
         Mult_Buf[14].Feature_n = FeatureBuf_602;
         Mult_Buf[14].Weight_n = Wgt_4_602;
         Mult_Buf[15].Feature_n = FeatureBuf_603;
         Mult_Buf[15].Weight_n = Wgt_4_603;
         Mult_Buf[16].Feature_n = FeatureBuf_604;
         Mult_Buf[16].Weight_n = Wgt_4_604;
         Mult_Buf[17].Feature_n = FeatureBuf_605;
         Mult_Buf[17].Weight_n = Wgt_4_605;
         Mult_Buf[18].Feature_n = FeatureBuf_606;
         Mult_Buf[18].Weight_n = Wgt_4_606;
         Mult_Buf[19].Feature_n = FeatureBuf_607;
         Mult_Buf[19].Weight_n = Wgt_4_607;
         Mult_Buf[20].Feature_n = FeatureBuf_608;
         Mult_Buf[20].Weight_n = Wgt_4_608;
         Mult_Buf[21].Feature_n = FeatureBuf_609;
         Mult_Buf[21].Weight_n = Wgt_4_609;
         Mult_Buf[22].Feature_n = FeatureBuf_610;
         Mult_Buf[22].Weight_n = Wgt_4_610;
         Mult_Buf[23].Feature_n = FeatureBuf_611;
         Mult_Buf[23].Weight_n = Wgt_4_611;
         Mult_Buf[24].Feature_n = FeatureBuf_612;
         Mult_Buf[24].Weight_n = Wgt_4_612;
         Mult_Buf[25].Feature_n = FeatureBuf_613;
         Mult_Buf[25].Weight_n = Wgt_4_613;
         Mult_Buf[26].Feature_n = FeatureBuf_614;
         Mult_Buf[26].Weight_n = Wgt_4_614;
         Mult_Buf[27].Feature_n = FeatureBuf_615;
         Mult_Buf[27].Weight_n = Wgt_4_615;
         Mult_Buf[28].Feature_n = FeatureBuf_616;
         Mult_Buf[28].Weight_n = Wgt_4_616;
         Mult_Buf[29].Feature_n = FeatureBuf_617;
         Mult_Buf[29].Weight_n = Wgt_4_617;
         Mult_Buf[30].Feature_n = FeatureBuf_618;
         Mult_Buf[30].Weight_n = Wgt_4_618;
         Mult_Buf[31].Feature_n = FeatureBuf_619;
         Mult_Buf[31].Weight_n = Wgt_4_619;
         Mult_Buf[32].Feature_n = FeatureBuf_620;
         Mult_Buf[32].Weight_n = Wgt_4_620;
         Mult_Buf[33].Feature_n = FeatureBuf_621;
         Mult_Buf[33].Weight_n = Wgt_4_621;
         Mult_Buf[34].Feature_n = FeatureBuf_622;
         Mult_Buf[34].Weight_n = Wgt_4_622;
         Mult_Buf[35].Feature_n = FeatureBuf_623;
         Mult_Buf[35].Weight_n = Wgt_4_623;
         Mult_Buf[36].Feature_n = FeatureBuf_624;
         Mult_Buf[36].Weight_n = Wgt_4_624;
         Mult_Buf[37].Feature_n = FeatureBuf_625;
         Mult_Buf[37].Weight_n = Wgt_4_625;
         Mult_Buf[38].Feature_n = FeatureBuf_626;
         Mult_Buf[38].Weight_n = Wgt_4_626;
         Mult_Buf[39].Feature_n = FeatureBuf_627;
         Mult_Buf[39].Weight_n = Wgt_4_627;
         Mult_Buf[40].Feature_n = FeatureBuf_628;
         Mult_Buf[40].Weight_n = Wgt_4_628;
         Mult_Buf[41].Feature_n = FeatureBuf_629;
         Mult_Buf[41].Weight_n = Wgt_4_629;
         Mult_Buf[42].Feature_n = FeatureBuf_630;
         Mult_Buf[42].Weight_n = Wgt_4_630;
         Mult_Buf[43].Feature_n = FeatureBuf_631;
         Mult_Buf[43].Weight_n = Wgt_4_631;
         Mult_Buf[44].Feature_n = FeatureBuf_632;
         Mult_Buf[44].Weight_n = Wgt_4_632;
         Mult_Buf[45].Feature_n = FeatureBuf_633;
         Mult_Buf[45].Weight_n = Wgt_4_633;
         Mult_Buf[46].Feature_n = FeatureBuf_634;
         Mult_Buf[46].Weight_n = Wgt_4_634;
         Mult_Buf[47].Feature_n = FeatureBuf_635;
         Mult_Buf[47].Weight_n = Wgt_4_635;
         Mult_Buf[48].Feature_n = FeatureBuf_636;
         Mult_Buf[48].Weight_n = Wgt_4_636;
         Mult_Buf[49].Feature_n = FeatureBuf_637;
         Mult_Buf[49].Weight_n = Wgt_4_637;
         Mult_Buf[50].Feature_n = FeatureBuf_638;
         Mult_Buf[50].Weight_n = Wgt_4_638;
         Mult_Buf[51].Feature_n = FeatureBuf_639;
         Mult_Buf[51].Weight_n = Wgt_4_639;
         Mult_Buf[52].Feature_n = FeatureBuf_640;
         Mult_Buf[52].Weight_n = Wgt_4_640;
         Mult_Buf[53].Feature_n = FeatureBuf_641;
         Mult_Buf[53].Weight_n = Wgt_4_641;
         Mult_Buf[54].Feature_n = FeatureBuf_642;
         Mult_Buf[54].Weight_n = Wgt_4_642;
         Mult_Buf[55].Feature_n = FeatureBuf_643;
         Mult_Buf[55].Weight_n = Wgt_4_643;
         Mult_Buf[56].Feature_n = FeatureBuf_644;
         Mult_Buf[56].Weight_n = Wgt_4_644;
         Mult_Buf[57].Feature_n = FeatureBuf_645;
         Mult_Buf[57].Weight_n = Wgt_4_645;
         Mult_Buf[58].Feature_n = FeatureBuf_646;
         Mult_Buf[58].Weight_n = Wgt_4_646;
         Mult_Buf[59].Feature_n = FeatureBuf_647;
         Mult_Buf[59].Weight_n = Wgt_4_647;
         Mult_Buf[60].Feature_n = FeatureBuf_648;
         Mult_Buf[60].Weight_n = Wgt_4_648;
         Mult_Buf[61].Feature_n = FeatureBuf_649;
         Mult_Buf[61].Weight_n = Wgt_4_649;
         Mult_Buf[62].Feature_n = FeatureBuf_650;
         Mult_Buf[62].Weight_n = Wgt_4_650;
         Mult_Buf[63].Feature_n = FeatureBuf_651;
         Mult_Buf[63].Weight_n = Wgt_4_651;
         Mult_Buf[64].Feature_n = FeatureBuf_652;
         Mult_Buf[64].Weight_n = Wgt_4_652;
         Mult_Buf[65].Feature_n = FeatureBuf_653;
         Mult_Buf[65].Weight_n = Wgt_4_653;
         Mult_Buf[66].Feature_n = FeatureBuf_654;
         Mult_Buf[66].Weight_n = Wgt_4_654;
         Mult_Buf[67].Feature_n = FeatureBuf_655;
         Mult_Buf[67].Weight_n = Wgt_4_655;
         Mult_Buf[68].Feature_n = FeatureBuf_656;
         Mult_Buf[68].Weight_n = Wgt_4_656;
         Mult_Buf[69].Feature_n = FeatureBuf_657;
         Mult_Buf[69].Weight_n = Wgt_4_657;
         Mult_Buf[70].Feature_n = FeatureBuf_658;
         Mult_Buf[70].Weight_n = Wgt_4_658;
         Mult_Buf[71].Feature_n = FeatureBuf_659;
         Mult_Buf[71].Weight_n = Wgt_4_659;
         Mult_Buf[72].Feature_n = FeatureBuf_660;
         Mult_Buf[72].Weight_n = Wgt_4_660;
         Mult_Buf[73].Feature_n = FeatureBuf_661;
         Mult_Buf[73].Weight_n = Wgt_4_661;
         Mult_Buf[74].Feature_n = FeatureBuf_662;
         Mult_Buf[74].Weight_n = Wgt_4_662;
         Mult_Buf[75].Feature_n = FeatureBuf_663;
         Mult_Buf[75].Weight_n = Wgt_4_663;
         Mult_Buf[76].Feature_n = FeatureBuf_664;
         Mult_Buf[76].Weight_n = Wgt_4_664;
         Mult_Buf[77].Feature_n = FeatureBuf_665;
         Mult_Buf[77].Weight_n = Wgt_4_665;
         Mult_Buf[78].Feature_n = FeatureBuf_666;
         Mult_Buf[78].Weight_n = Wgt_4_666;
         Mult_Buf[79].Feature_n = FeatureBuf_667;
         Mult_Buf[79].Weight_n = Wgt_4_667;
         Mult_Buf[80].Feature_n = FeatureBuf_668;
         Mult_Buf[80].Weight_n = Wgt_4_668;
         Mult_Buf[81].Feature_n = FeatureBuf_669;
         Mult_Buf[81].Weight_n = Wgt_4_669;
         Mult_Buf[82].Feature_n = FeatureBuf_670;
         Mult_Buf[82].Weight_n = Wgt_4_670;
         Mult_Buf[83].Feature_n = FeatureBuf_671;
         Mult_Buf[83].Weight_n = Wgt_4_671;
         Mult_Buf[84].Feature_n = FeatureBuf_672;
         Mult_Buf[84].Weight_n = Wgt_4_672;
         Mult_Buf[85].Feature_n = FeatureBuf_673;
         Mult_Buf[85].Weight_n = Wgt_4_673;
         Mult_Buf[86].Feature_n = FeatureBuf_674;
         Mult_Buf[86].Weight_n = Wgt_4_674;
         Mult_Buf[87].Feature_n = FeatureBuf_675;
         Mult_Buf[87].Weight_n = Wgt_4_675;
         Mult_Buf[88].Feature_n = FeatureBuf_676;
         Mult_Buf[88].Weight_n = Wgt_4_676;
         Mult_Buf[89].Feature_n = FeatureBuf_677;
         Mult_Buf[89].Weight_n = Wgt_4_677;
         Mult_Buf[90].Feature_n = FeatureBuf_678;
         Mult_Buf[90].Weight_n = Wgt_4_678;
         Mult_Buf[91].Feature_n = FeatureBuf_679;
         Mult_Buf[91].Weight_n = Wgt_4_679;
         Mult_Buf[92].Feature_n = FeatureBuf_680;
         Mult_Buf[92].Weight_n = Wgt_4_680;
         Mult_Buf[93].Feature_n = FeatureBuf_681;
         Mult_Buf[93].Weight_n = Wgt_4_681;
         Mult_Buf[94].Feature_n = FeatureBuf_682;
         Mult_Buf[94].Weight_n = Wgt_4_682;
         Mult_Buf[95].Feature_n = FeatureBuf_683;
         Mult_Buf[95].Weight_n = Wgt_4_683;
         Mult_Buf[96].Feature_n = FeatureBuf_684;
         Mult_Buf[96].Weight_n = Wgt_4_684;
         Mult_Buf[97].Feature_n = FeatureBuf_685;
         Mult_Buf[97].Weight_n = Wgt_4_685;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     //Collect Partial result form Adder
         Res_2_0_n = Part_Res;
     end
    41:begin
     nxt_state = 42;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_686;
         Mult_Buf[0].Weight_n = Wgt_4_686;
         Mult_Buf[1].Feature_n = FeatureBuf_687;
         Mult_Buf[1].Weight_n = Wgt_4_687;
         Mult_Buf[2].Feature_n = FeatureBuf_688;
         Mult_Buf[2].Weight_n = Wgt_4_688;
         Mult_Buf[3].Feature_n = FeatureBuf_689;
         Mult_Buf[3].Weight_n = Wgt_4_689;
         Mult_Buf[4].Feature_n = FeatureBuf_690;
         Mult_Buf[4].Weight_n = Wgt_4_690;
         Mult_Buf[5].Feature_n = FeatureBuf_691;
         Mult_Buf[5].Weight_n = Wgt_4_691;
         Mult_Buf[6].Feature_n = FeatureBuf_692;
         Mult_Buf[6].Weight_n = Wgt_4_692;
         Mult_Buf[7].Feature_n = FeatureBuf_693;
         Mult_Buf[7].Weight_n = Wgt_4_693;
         Mult_Buf[8].Feature_n = FeatureBuf_694;
         Mult_Buf[8].Weight_n = Wgt_4_694;
         Mult_Buf[9].Feature_n = FeatureBuf_695;
         Mult_Buf[9].Weight_n = Wgt_4_695;
         Mult_Buf[10].Feature_n = FeatureBuf_696;
         Mult_Buf[10].Weight_n = Wgt_4_696;
         Mult_Buf[11].Feature_n = FeatureBuf_697;
         Mult_Buf[11].Weight_n = Wgt_4_697;
         Mult_Buf[12].Feature_n = FeatureBuf_698;
         Mult_Buf[12].Weight_n = Wgt_4_698;
         Mult_Buf[13].Feature_n = FeatureBuf_699;
         Mult_Buf[13].Weight_n = Wgt_4_699;
         Mult_Buf[14].Feature_n = FeatureBuf_700;
         Mult_Buf[14].Weight_n = Wgt_4_700;
         Mult_Buf[15].Feature_n = FeatureBuf_701;
         Mult_Buf[15].Weight_n = Wgt_4_701;
         Mult_Buf[16].Feature_n = FeatureBuf_702;
         Mult_Buf[16].Weight_n = Wgt_4_702;
         Mult_Buf[17].Feature_n = FeatureBuf_703;
         Mult_Buf[17].Weight_n = Wgt_4_703;
         Mult_Buf[18].Feature_n = FeatureBuf_704;
         Mult_Buf[18].Weight_n = Wgt_4_704;
         Mult_Buf[19].Feature_n = FeatureBuf_705;
         Mult_Buf[19].Weight_n = Wgt_4_705;
         Mult_Buf[20].Feature_n = FeatureBuf_706;
         Mult_Buf[20].Weight_n = Wgt_4_706;
         Mult_Buf[21].Feature_n = FeatureBuf_707;
         Mult_Buf[21].Weight_n = Wgt_4_707;
         Mult_Buf[22].Feature_n = FeatureBuf_708;
         Mult_Buf[22].Weight_n = Wgt_4_708;
         Mult_Buf[23].Feature_n = FeatureBuf_709;
         Mult_Buf[23].Weight_n = Wgt_4_709;
         Mult_Buf[24].Feature_n = FeatureBuf_710;
         Mult_Buf[24].Weight_n = Wgt_4_710;
         Mult_Buf[25].Feature_n = FeatureBuf_711;
         Mult_Buf[25].Weight_n = Wgt_4_711;
         Mult_Buf[26].Feature_n = FeatureBuf_712;
         Mult_Buf[26].Weight_n = Wgt_4_712;
         Mult_Buf[27].Feature_n = FeatureBuf_713;
         Mult_Buf[27].Weight_n = Wgt_4_713;
         Mult_Buf[28].Feature_n = FeatureBuf_714;
         Mult_Buf[28].Weight_n = Wgt_4_714;
         Mult_Buf[29].Feature_n = FeatureBuf_715;
         Mult_Buf[29].Weight_n = Wgt_4_715;
         Mult_Buf[30].Feature_n = FeatureBuf_716;
         Mult_Buf[30].Weight_n = Wgt_4_716;
         Mult_Buf[31].Feature_n = FeatureBuf_717;
         Mult_Buf[31].Weight_n = Wgt_4_717;
         Mult_Buf[32].Feature_n = FeatureBuf_718;
         Mult_Buf[32].Weight_n = Wgt_4_718;
         Mult_Buf[33].Feature_n = FeatureBuf_719;
         Mult_Buf[33].Weight_n = Wgt_4_719;
         Mult_Buf[34].Feature_n = FeatureBuf_720;
         Mult_Buf[34].Weight_n = Wgt_4_720;
         Mult_Buf[35].Feature_n = FeatureBuf_721;
         Mult_Buf[35].Weight_n = Wgt_4_721;
         Mult_Buf[36].Feature_n = FeatureBuf_722;
         Mult_Buf[36].Weight_n = Wgt_4_722;
         Mult_Buf[37].Feature_n = FeatureBuf_723;
         Mult_Buf[37].Weight_n = Wgt_4_723;
         Mult_Buf[38].Feature_n = FeatureBuf_724;
         Mult_Buf[38].Weight_n = Wgt_4_724;
         Mult_Buf[39].Feature_n = FeatureBuf_725;
         Mult_Buf[39].Weight_n = Wgt_4_725;
         Mult_Buf[40].Feature_n = FeatureBuf_726;
         Mult_Buf[40].Weight_n = Wgt_4_726;
         Mult_Buf[41].Feature_n = FeatureBuf_727;
         Mult_Buf[41].Weight_n = Wgt_4_727;
         Mult_Buf[42].Feature_n = FeatureBuf_728;
         Mult_Buf[42].Weight_n = Wgt_4_728;
         Mult_Buf[43].Feature_n = FeatureBuf_729;
         Mult_Buf[43].Weight_n = Wgt_4_729;
         Mult_Buf[44].Feature_n = FeatureBuf_730;
         Mult_Buf[44].Weight_n = Wgt_4_730;
         Mult_Buf[45].Feature_n = FeatureBuf_731;
         Mult_Buf[45].Weight_n = Wgt_4_731;
         Mult_Buf[46].Feature_n = FeatureBuf_732;
         Mult_Buf[46].Weight_n = Wgt_4_732;
         Mult_Buf[47].Feature_n = FeatureBuf_733;
         Mult_Buf[47].Weight_n = Wgt_4_733;
         Mult_Buf[48].Feature_n = FeatureBuf_734;
         Mult_Buf[48].Weight_n = Wgt_4_734;
         Mult_Buf[49].Feature_n = FeatureBuf_735;
         Mult_Buf[49].Weight_n = Wgt_4_735;
         Mult_Buf[50].Feature_n = FeatureBuf_736;
         Mult_Buf[50].Weight_n = Wgt_4_736;
         Mult_Buf[51].Feature_n = FeatureBuf_737;
         Mult_Buf[51].Weight_n = Wgt_4_737;
         Mult_Buf[52].Feature_n = FeatureBuf_738;
         Mult_Buf[52].Weight_n = Wgt_4_738;
         Mult_Buf[53].Feature_n = FeatureBuf_739;
         Mult_Buf[53].Weight_n = Wgt_4_739;
         Mult_Buf[54].Feature_n = FeatureBuf_740;
         Mult_Buf[54].Weight_n = Wgt_4_740;
         Mult_Buf[55].Feature_n = FeatureBuf_741;
         Mult_Buf[55].Weight_n = Wgt_4_741;
         Mult_Buf[56].Feature_n = FeatureBuf_742;
         Mult_Buf[56].Weight_n = Wgt_4_742;
         Mult_Buf[57].Feature_n = FeatureBuf_743;
         Mult_Buf[57].Weight_n = Wgt_4_743;
         Mult_Buf[58].Feature_n = FeatureBuf_744;
         Mult_Buf[58].Weight_n = Wgt_4_744;
         Mult_Buf[59].Feature_n = FeatureBuf_745;
         Mult_Buf[59].Weight_n = Wgt_4_745;
         Mult_Buf[60].Feature_n = FeatureBuf_746;
         Mult_Buf[60].Weight_n = Wgt_4_746;
         Mult_Buf[61].Feature_n = FeatureBuf_747;
         Mult_Buf[61].Weight_n = Wgt_4_747;
         Mult_Buf[62].Feature_n = FeatureBuf_748;
         Mult_Buf[62].Weight_n = Wgt_4_748;
         Mult_Buf[63].Feature_n = FeatureBuf_749;
         Mult_Buf[63].Weight_n = Wgt_4_749;
         Mult_Buf[64].Feature_n = FeatureBuf_750;
         Mult_Buf[64].Weight_n = Wgt_4_750;
         Mult_Buf[65].Feature_n = FeatureBuf_751;
         Mult_Buf[65].Weight_n = Wgt_4_751;
         Mult_Buf[66].Feature_n = FeatureBuf_752;
         Mult_Buf[66].Weight_n = Wgt_4_752;
         Mult_Buf[67].Feature_n = FeatureBuf_753;
         Mult_Buf[67].Weight_n = Wgt_4_753;
         Mult_Buf[68].Feature_n = FeatureBuf_754;
         Mult_Buf[68].Weight_n = Wgt_4_754;
         Mult_Buf[69].Feature_n = FeatureBuf_755;
         Mult_Buf[69].Weight_n = Wgt_4_755;
         Mult_Buf[70].Feature_n = FeatureBuf_756;
         Mult_Buf[70].Weight_n = Wgt_4_756;
         Mult_Buf[71].Feature_n = FeatureBuf_757;
         Mult_Buf[71].Weight_n = Wgt_4_757;
         Mult_Buf[72].Feature_n = FeatureBuf_758;
         Mult_Buf[72].Weight_n = Wgt_4_758;
         Mult_Buf[73].Feature_n = FeatureBuf_759;
         Mult_Buf[73].Weight_n = Wgt_4_759;
         Mult_Buf[74].Feature_n = FeatureBuf_760;
         Mult_Buf[74].Weight_n = Wgt_4_760;
         Mult_Buf[75].Feature_n = FeatureBuf_761;
         Mult_Buf[75].Weight_n = Wgt_4_761;
         Mult_Buf[76].Feature_n = FeatureBuf_762;
         Mult_Buf[76].Weight_n = Wgt_4_762;
         Mult_Buf[77].Feature_n = FeatureBuf_763;
         Mult_Buf[77].Weight_n = Wgt_4_763;
         Mult_Buf[78].Feature_n = FeatureBuf_764;
         Mult_Buf[78].Weight_n = Wgt_4_764;
         Mult_Buf[79].Feature_n = FeatureBuf_765;
         Mult_Buf[79].Weight_n = Wgt_4_765;
         Mult_Buf[80].Feature_n = FeatureBuf_766;
         Mult_Buf[80].Weight_n = Wgt_4_766;
         Mult_Buf[81].Feature_n = FeatureBuf_767;
         Mult_Buf[81].Weight_n = Wgt_4_767;
         Mult_Buf[82].Feature_n = FeatureBuf_768;
         Mult_Buf[82].Weight_n = Wgt_4_768;
         Mult_Buf[83].Feature_n = FeatureBuf_769;
         Mult_Buf[83].Weight_n = Wgt_4_769;
         Mult_Buf[84].Feature_n = FeatureBuf_770;
         Mult_Buf[84].Weight_n = Wgt_4_770;
         Mult_Buf[85].Feature_n = FeatureBuf_771;
         Mult_Buf[85].Weight_n = Wgt_4_771;
         Mult_Buf[86].Feature_n = FeatureBuf_772;
         Mult_Buf[86].Weight_n = Wgt_4_772;
         Mult_Buf[87].Feature_n = FeatureBuf_773;
         Mult_Buf[87].Weight_n = Wgt_4_773;
         Mult_Buf[88].Feature_n = FeatureBuf_774;
         Mult_Buf[88].Weight_n = Wgt_4_774;
         Mult_Buf[89].Feature_n = FeatureBuf_775;
         Mult_Buf[89].Weight_n = Wgt_4_775;
         Mult_Buf[90].Feature_n = FeatureBuf_776;
         Mult_Buf[90].Weight_n = Wgt_4_776;
         Mult_Buf[91].Feature_n = FeatureBuf_777;
         Mult_Buf[91].Weight_n = Wgt_4_777;
         Mult_Buf[92].Feature_n = FeatureBuf_778;
         Mult_Buf[92].Weight_n = Wgt_4_778;
         Mult_Buf[93].Feature_n = FeatureBuf_779;
         Mult_Buf[93].Weight_n = Wgt_4_779;
         Mult_Buf[94].Feature_n = FeatureBuf_780;
         Mult_Buf[94].Weight_n = Wgt_4_780;
         Mult_Buf[95].Feature_n = FeatureBuf_781;
         Mult_Buf[95].Weight_n = Wgt_4_781;
         Mult_Buf[96].Feature_n = FeatureBuf_782;
         Mult_Buf[96].Weight_n = Wgt_4_782;
         Mult_Buf[97].Feature_n = FeatureBuf_783;
         Mult_Buf[97].Weight_n = Wgt_4_783;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     //Collect Partial result form Adder
         Res_2_1_n = Part_Res;
     end
    42:begin
     nxt_state = 43;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_0;
         Mult_Buf[0].Weight_n = Wgt_5_0;
         Mult_Buf[1].Feature_n = FeatureBuf_1;
         Mult_Buf[1].Weight_n = Wgt_5_1;
         Mult_Buf[2].Feature_n = FeatureBuf_2;
         Mult_Buf[2].Weight_n = Wgt_5_2;
         Mult_Buf[3].Feature_n = FeatureBuf_3;
         Mult_Buf[3].Weight_n = Wgt_5_3;
         Mult_Buf[4].Feature_n = FeatureBuf_4;
         Mult_Buf[4].Weight_n = Wgt_5_4;
         Mult_Buf[5].Feature_n = FeatureBuf_5;
         Mult_Buf[5].Weight_n = Wgt_5_5;
         Mult_Buf[6].Feature_n = FeatureBuf_6;
         Mult_Buf[6].Weight_n = Wgt_5_6;
         Mult_Buf[7].Feature_n = FeatureBuf_7;
         Mult_Buf[7].Weight_n = Wgt_5_7;
         Mult_Buf[8].Feature_n = FeatureBuf_8;
         Mult_Buf[8].Weight_n = Wgt_5_8;
         Mult_Buf[9].Feature_n = FeatureBuf_9;
         Mult_Buf[9].Weight_n = Wgt_5_9;
         Mult_Buf[10].Feature_n = FeatureBuf_10;
         Mult_Buf[10].Weight_n = Wgt_5_10;
         Mult_Buf[11].Feature_n = FeatureBuf_11;
         Mult_Buf[11].Weight_n = Wgt_5_11;
         Mult_Buf[12].Feature_n = FeatureBuf_12;
         Mult_Buf[12].Weight_n = Wgt_5_12;
         Mult_Buf[13].Feature_n = FeatureBuf_13;
         Mult_Buf[13].Weight_n = Wgt_5_13;
         Mult_Buf[14].Feature_n = FeatureBuf_14;
         Mult_Buf[14].Weight_n = Wgt_5_14;
         Mult_Buf[15].Feature_n = FeatureBuf_15;
         Mult_Buf[15].Weight_n = Wgt_5_15;
         Mult_Buf[16].Feature_n = FeatureBuf_16;
         Mult_Buf[16].Weight_n = Wgt_5_16;
         Mult_Buf[17].Feature_n = FeatureBuf_17;
         Mult_Buf[17].Weight_n = Wgt_5_17;
         Mult_Buf[18].Feature_n = FeatureBuf_18;
         Mult_Buf[18].Weight_n = Wgt_5_18;
         Mult_Buf[19].Feature_n = FeatureBuf_19;
         Mult_Buf[19].Weight_n = Wgt_5_19;
         Mult_Buf[20].Feature_n = FeatureBuf_20;
         Mult_Buf[20].Weight_n = Wgt_5_20;
         Mult_Buf[21].Feature_n = FeatureBuf_21;
         Mult_Buf[21].Weight_n = Wgt_5_21;
         Mult_Buf[22].Feature_n = FeatureBuf_22;
         Mult_Buf[22].Weight_n = Wgt_5_22;
         Mult_Buf[23].Feature_n = FeatureBuf_23;
         Mult_Buf[23].Weight_n = Wgt_5_23;
         Mult_Buf[24].Feature_n = FeatureBuf_24;
         Mult_Buf[24].Weight_n = Wgt_5_24;
         Mult_Buf[25].Feature_n = FeatureBuf_25;
         Mult_Buf[25].Weight_n = Wgt_5_25;
         Mult_Buf[26].Feature_n = FeatureBuf_26;
         Mult_Buf[26].Weight_n = Wgt_5_26;
         Mult_Buf[27].Feature_n = FeatureBuf_27;
         Mult_Buf[27].Weight_n = Wgt_5_27;
         Mult_Buf[28].Feature_n = FeatureBuf_28;
         Mult_Buf[28].Weight_n = Wgt_5_28;
         Mult_Buf[29].Feature_n = FeatureBuf_29;
         Mult_Buf[29].Weight_n = Wgt_5_29;
         Mult_Buf[30].Feature_n = FeatureBuf_30;
         Mult_Buf[30].Weight_n = Wgt_5_30;
         Mult_Buf[31].Feature_n = FeatureBuf_31;
         Mult_Buf[31].Weight_n = Wgt_5_31;
         Mult_Buf[32].Feature_n = FeatureBuf_32;
         Mult_Buf[32].Weight_n = Wgt_5_32;
         Mult_Buf[33].Feature_n = FeatureBuf_33;
         Mult_Buf[33].Weight_n = Wgt_5_33;
         Mult_Buf[34].Feature_n = FeatureBuf_34;
         Mult_Buf[34].Weight_n = Wgt_5_34;
         Mult_Buf[35].Feature_n = FeatureBuf_35;
         Mult_Buf[35].Weight_n = Wgt_5_35;
         Mult_Buf[36].Feature_n = FeatureBuf_36;
         Mult_Buf[36].Weight_n = Wgt_5_36;
         Mult_Buf[37].Feature_n = FeatureBuf_37;
         Mult_Buf[37].Weight_n = Wgt_5_37;
         Mult_Buf[38].Feature_n = FeatureBuf_38;
         Mult_Buf[38].Weight_n = Wgt_5_38;
         Mult_Buf[39].Feature_n = FeatureBuf_39;
         Mult_Buf[39].Weight_n = Wgt_5_39;
         Mult_Buf[40].Feature_n = FeatureBuf_40;
         Mult_Buf[40].Weight_n = Wgt_5_40;
         Mult_Buf[41].Feature_n = FeatureBuf_41;
         Mult_Buf[41].Weight_n = Wgt_5_41;
         Mult_Buf[42].Feature_n = FeatureBuf_42;
         Mult_Buf[42].Weight_n = Wgt_5_42;
         Mult_Buf[43].Feature_n = FeatureBuf_43;
         Mult_Buf[43].Weight_n = Wgt_5_43;
         Mult_Buf[44].Feature_n = FeatureBuf_44;
         Mult_Buf[44].Weight_n = Wgt_5_44;
         Mult_Buf[45].Feature_n = FeatureBuf_45;
         Mult_Buf[45].Weight_n = Wgt_5_45;
         Mult_Buf[46].Feature_n = FeatureBuf_46;
         Mult_Buf[46].Weight_n = Wgt_5_46;
         Mult_Buf[47].Feature_n = FeatureBuf_47;
         Mult_Buf[47].Weight_n = Wgt_5_47;
         Mult_Buf[48].Feature_n = FeatureBuf_48;
         Mult_Buf[48].Weight_n = Wgt_5_48;
         Mult_Buf[49].Feature_n = FeatureBuf_49;
         Mult_Buf[49].Weight_n = Wgt_5_49;
         Mult_Buf[50].Feature_n = FeatureBuf_50;
         Mult_Buf[50].Weight_n = Wgt_5_50;
         Mult_Buf[51].Feature_n = FeatureBuf_51;
         Mult_Buf[51].Weight_n = Wgt_5_51;
         Mult_Buf[52].Feature_n = FeatureBuf_52;
         Mult_Buf[52].Weight_n = Wgt_5_52;
         Mult_Buf[53].Feature_n = FeatureBuf_53;
         Mult_Buf[53].Weight_n = Wgt_5_53;
         Mult_Buf[54].Feature_n = FeatureBuf_54;
         Mult_Buf[54].Weight_n = Wgt_5_54;
         Mult_Buf[55].Feature_n = FeatureBuf_55;
         Mult_Buf[55].Weight_n = Wgt_5_55;
         Mult_Buf[56].Feature_n = FeatureBuf_56;
         Mult_Buf[56].Weight_n = Wgt_5_56;
         Mult_Buf[57].Feature_n = FeatureBuf_57;
         Mult_Buf[57].Weight_n = Wgt_5_57;
         Mult_Buf[58].Feature_n = FeatureBuf_58;
         Mult_Buf[58].Weight_n = Wgt_5_58;
         Mult_Buf[59].Feature_n = FeatureBuf_59;
         Mult_Buf[59].Weight_n = Wgt_5_59;
         Mult_Buf[60].Feature_n = FeatureBuf_60;
         Mult_Buf[60].Weight_n = Wgt_5_60;
         Mult_Buf[61].Feature_n = FeatureBuf_61;
         Mult_Buf[61].Weight_n = Wgt_5_61;
         Mult_Buf[62].Feature_n = FeatureBuf_62;
         Mult_Buf[62].Weight_n = Wgt_5_62;
         Mult_Buf[63].Feature_n = FeatureBuf_63;
         Mult_Buf[63].Weight_n = Wgt_5_63;
         Mult_Buf[64].Feature_n = FeatureBuf_64;
         Mult_Buf[64].Weight_n = Wgt_5_64;
         Mult_Buf[65].Feature_n = FeatureBuf_65;
         Mult_Buf[65].Weight_n = Wgt_5_65;
         Mult_Buf[66].Feature_n = FeatureBuf_66;
         Mult_Buf[66].Weight_n = Wgt_5_66;
         Mult_Buf[67].Feature_n = FeatureBuf_67;
         Mult_Buf[67].Weight_n = Wgt_5_67;
         Mult_Buf[68].Feature_n = FeatureBuf_68;
         Mult_Buf[68].Weight_n = Wgt_5_68;
         Mult_Buf[69].Feature_n = FeatureBuf_69;
         Mult_Buf[69].Weight_n = Wgt_5_69;
         Mult_Buf[70].Feature_n = FeatureBuf_70;
         Mult_Buf[70].Weight_n = Wgt_5_70;
         Mult_Buf[71].Feature_n = FeatureBuf_71;
         Mult_Buf[71].Weight_n = Wgt_5_71;
         Mult_Buf[72].Feature_n = FeatureBuf_72;
         Mult_Buf[72].Weight_n = Wgt_5_72;
         Mult_Buf[73].Feature_n = FeatureBuf_73;
         Mult_Buf[73].Weight_n = Wgt_5_73;
         Mult_Buf[74].Feature_n = FeatureBuf_74;
         Mult_Buf[74].Weight_n = Wgt_5_74;
         Mult_Buf[75].Feature_n = FeatureBuf_75;
         Mult_Buf[75].Weight_n = Wgt_5_75;
         Mult_Buf[76].Feature_n = FeatureBuf_76;
         Mult_Buf[76].Weight_n = Wgt_5_76;
         Mult_Buf[77].Feature_n = FeatureBuf_77;
         Mult_Buf[77].Weight_n = Wgt_5_77;
         Mult_Buf[78].Feature_n = FeatureBuf_78;
         Mult_Buf[78].Weight_n = Wgt_5_78;
         Mult_Buf[79].Feature_n = FeatureBuf_79;
         Mult_Buf[79].Weight_n = Wgt_5_79;
         Mult_Buf[80].Feature_n = FeatureBuf_80;
         Mult_Buf[80].Weight_n = Wgt_5_80;
         Mult_Buf[81].Feature_n = FeatureBuf_81;
         Mult_Buf[81].Weight_n = Wgt_5_81;
         Mult_Buf[82].Feature_n = FeatureBuf_82;
         Mult_Buf[82].Weight_n = Wgt_5_82;
         Mult_Buf[83].Feature_n = FeatureBuf_83;
         Mult_Buf[83].Weight_n = Wgt_5_83;
         Mult_Buf[84].Feature_n = FeatureBuf_84;
         Mult_Buf[84].Weight_n = Wgt_5_84;
         Mult_Buf[85].Feature_n = FeatureBuf_85;
         Mult_Buf[85].Weight_n = Wgt_5_85;
         Mult_Buf[86].Feature_n = FeatureBuf_86;
         Mult_Buf[86].Weight_n = Wgt_5_86;
         Mult_Buf[87].Feature_n = FeatureBuf_87;
         Mult_Buf[87].Weight_n = Wgt_5_87;
         Mult_Buf[88].Feature_n = FeatureBuf_88;
         Mult_Buf[88].Weight_n = Wgt_5_88;
         Mult_Buf[89].Feature_n = FeatureBuf_89;
         Mult_Buf[89].Weight_n = Wgt_5_89;
         Mult_Buf[90].Feature_n = FeatureBuf_90;
         Mult_Buf[90].Weight_n = Wgt_5_90;
         Mult_Buf[91].Feature_n = FeatureBuf_91;
         Mult_Buf[91].Weight_n = Wgt_5_91;
         Mult_Buf[92].Feature_n = FeatureBuf_92;
         Mult_Buf[92].Weight_n = Wgt_5_92;
         Mult_Buf[93].Feature_n = FeatureBuf_93;
         Mult_Buf[93].Weight_n = Wgt_5_93;
         Mult_Buf[94].Feature_n = FeatureBuf_94;
         Mult_Buf[94].Weight_n = Wgt_5_94;
         Mult_Buf[95].Feature_n = FeatureBuf_95;
         Mult_Buf[95].Weight_n = Wgt_5_95;
         Mult_Buf[96].Feature_n = FeatureBuf_96;
         Mult_Buf[96].Weight_n = Wgt_5_96;
         Mult_Buf[97].Feature_n = FeatureBuf_97;
         Mult_Buf[97].Weight_n = Wgt_5_97;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     //Collect Partial result form Adder
         Res_2_2_n = Part_Res;
     end
    43:begin
     nxt_state = 44;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_98;
         Mult_Buf[0].Weight_n = Wgt_5_98;
         Mult_Buf[1].Feature_n = FeatureBuf_99;
         Mult_Buf[1].Weight_n = Wgt_5_99;
         Mult_Buf[2].Feature_n = FeatureBuf_100;
         Mult_Buf[2].Weight_n = Wgt_5_100;
         Mult_Buf[3].Feature_n = FeatureBuf_101;
         Mult_Buf[3].Weight_n = Wgt_5_101;
         Mult_Buf[4].Feature_n = FeatureBuf_102;
         Mult_Buf[4].Weight_n = Wgt_5_102;
         Mult_Buf[5].Feature_n = FeatureBuf_103;
         Mult_Buf[5].Weight_n = Wgt_5_103;
         Mult_Buf[6].Feature_n = FeatureBuf_104;
         Mult_Buf[6].Weight_n = Wgt_5_104;
         Mult_Buf[7].Feature_n = FeatureBuf_105;
         Mult_Buf[7].Weight_n = Wgt_5_105;
         Mult_Buf[8].Feature_n = FeatureBuf_106;
         Mult_Buf[8].Weight_n = Wgt_5_106;
         Mult_Buf[9].Feature_n = FeatureBuf_107;
         Mult_Buf[9].Weight_n = Wgt_5_107;
         Mult_Buf[10].Feature_n = FeatureBuf_108;
         Mult_Buf[10].Weight_n = Wgt_5_108;
         Mult_Buf[11].Feature_n = FeatureBuf_109;
         Mult_Buf[11].Weight_n = Wgt_5_109;
         Mult_Buf[12].Feature_n = FeatureBuf_110;
         Mult_Buf[12].Weight_n = Wgt_5_110;
         Mult_Buf[13].Feature_n = FeatureBuf_111;
         Mult_Buf[13].Weight_n = Wgt_5_111;
         Mult_Buf[14].Feature_n = FeatureBuf_112;
         Mult_Buf[14].Weight_n = Wgt_5_112;
         Mult_Buf[15].Feature_n = FeatureBuf_113;
         Mult_Buf[15].Weight_n = Wgt_5_113;
         Mult_Buf[16].Feature_n = FeatureBuf_114;
         Mult_Buf[16].Weight_n = Wgt_5_114;
         Mult_Buf[17].Feature_n = FeatureBuf_115;
         Mult_Buf[17].Weight_n = Wgt_5_115;
         Mult_Buf[18].Feature_n = FeatureBuf_116;
         Mult_Buf[18].Weight_n = Wgt_5_116;
         Mult_Buf[19].Feature_n = FeatureBuf_117;
         Mult_Buf[19].Weight_n = Wgt_5_117;
         Mult_Buf[20].Feature_n = FeatureBuf_118;
         Mult_Buf[20].Weight_n = Wgt_5_118;
         Mult_Buf[21].Feature_n = FeatureBuf_119;
         Mult_Buf[21].Weight_n = Wgt_5_119;
         Mult_Buf[22].Feature_n = FeatureBuf_120;
         Mult_Buf[22].Weight_n = Wgt_5_120;
         Mult_Buf[23].Feature_n = FeatureBuf_121;
         Mult_Buf[23].Weight_n = Wgt_5_121;
         Mult_Buf[24].Feature_n = FeatureBuf_122;
         Mult_Buf[24].Weight_n = Wgt_5_122;
         Mult_Buf[25].Feature_n = FeatureBuf_123;
         Mult_Buf[25].Weight_n = Wgt_5_123;
         Mult_Buf[26].Feature_n = FeatureBuf_124;
         Mult_Buf[26].Weight_n = Wgt_5_124;
         Mult_Buf[27].Feature_n = FeatureBuf_125;
         Mult_Buf[27].Weight_n = Wgt_5_125;
         Mult_Buf[28].Feature_n = FeatureBuf_126;
         Mult_Buf[28].Weight_n = Wgt_5_126;
         Mult_Buf[29].Feature_n = FeatureBuf_127;
         Mult_Buf[29].Weight_n = Wgt_5_127;
         Mult_Buf[30].Feature_n = FeatureBuf_128;
         Mult_Buf[30].Weight_n = Wgt_5_128;
         Mult_Buf[31].Feature_n = FeatureBuf_129;
         Mult_Buf[31].Weight_n = Wgt_5_129;
         Mult_Buf[32].Feature_n = FeatureBuf_130;
         Mult_Buf[32].Weight_n = Wgt_5_130;
         Mult_Buf[33].Feature_n = FeatureBuf_131;
         Mult_Buf[33].Weight_n = Wgt_5_131;
         Mult_Buf[34].Feature_n = FeatureBuf_132;
         Mult_Buf[34].Weight_n = Wgt_5_132;
         Mult_Buf[35].Feature_n = FeatureBuf_133;
         Mult_Buf[35].Weight_n = Wgt_5_133;
         Mult_Buf[36].Feature_n = FeatureBuf_134;
         Mult_Buf[36].Weight_n = Wgt_5_134;
         Mult_Buf[37].Feature_n = FeatureBuf_135;
         Mult_Buf[37].Weight_n = Wgt_5_135;
         Mult_Buf[38].Feature_n = FeatureBuf_136;
         Mult_Buf[38].Weight_n = Wgt_5_136;
         Mult_Buf[39].Feature_n = FeatureBuf_137;
         Mult_Buf[39].Weight_n = Wgt_5_137;
         Mult_Buf[40].Feature_n = FeatureBuf_138;
         Mult_Buf[40].Weight_n = Wgt_5_138;
         Mult_Buf[41].Feature_n = FeatureBuf_139;
         Mult_Buf[41].Weight_n = Wgt_5_139;
         Mult_Buf[42].Feature_n = FeatureBuf_140;
         Mult_Buf[42].Weight_n = Wgt_5_140;
         Mult_Buf[43].Feature_n = FeatureBuf_141;
         Mult_Buf[43].Weight_n = Wgt_5_141;
         Mult_Buf[44].Feature_n = FeatureBuf_142;
         Mult_Buf[44].Weight_n = Wgt_5_142;
         Mult_Buf[45].Feature_n = FeatureBuf_143;
         Mult_Buf[45].Weight_n = Wgt_5_143;
         Mult_Buf[46].Feature_n = FeatureBuf_144;
         Mult_Buf[46].Weight_n = Wgt_5_144;
         Mult_Buf[47].Feature_n = FeatureBuf_145;
         Mult_Buf[47].Weight_n = Wgt_5_145;
         Mult_Buf[48].Feature_n = FeatureBuf_146;
         Mult_Buf[48].Weight_n = Wgt_5_146;
         Mult_Buf[49].Feature_n = FeatureBuf_147;
         Mult_Buf[49].Weight_n = Wgt_5_147;
         Mult_Buf[50].Feature_n = FeatureBuf_148;
         Mult_Buf[50].Weight_n = Wgt_5_148;
         Mult_Buf[51].Feature_n = FeatureBuf_149;
         Mult_Buf[51].Weight_n = Wgt_5_149;
         Mult_Buf[52].Feature_n = FeatureBuf_150;
         Mult_Buf[52].Weight_n = Wgt_5_150;
         Mult_Buf[53].Feature_n = FeatureBuf_151;
         Mult_Buf[53].Weight_n = Wgt_5_151;
         Mult_Buf[54].Feature_n = FeatureBuf_152;
         Mult_Buf[54].Weight_n = Wgt_5_152;
         Mult_Buf[55].Feature_n = FeatureBuf_153;
         Mult_Buf[55].Weight_n = Wgt_5_153;
         Mult_Buf[56].Feature_n = FeatureBuf_154;
         Mult_Buf[56].Weight_n = Wgt_5_154;
         Mult_Buf[57].Feature_n = FeatureBuf_155;
         Mult_Buf[57].Weight_n = Wgt_5_155;
         Mult_Buf[58].Feature_n = FeatureBuf_156;
         Mult_Buf[58].Weight_n = Wgt_5_156;
         Mult_Buf[59].Feature_n = FeatureBuf_157;
         Mult_Buf[59].Weight_n = Wgt_5_157;
         Mult_Buf[60].Feature_n = FeatureBuf_158;
         Mult_Buf[60].Weight_n = Wgt_5_158;
         Mult_Buf[61].Feature_n = FeatureBuf_159;
         Mult_Buf[61].Weight_n = Wgt_5_159;
         Mult_Buf[62].Feature_n = FeatureBuf_160;
         Mult_Buf[62].Weight_n = Wgt_5_160;
         Mult_Buf[63].Feature_n = FeatureBuf_161;
         Mult_Buf[63].Weight_n = Wgt_5_161;
         Mult_Buf[64].Feature_n = FeatureBuf_162;
         Mult_Buf[64].Weight_n = Wgt_5_162;
         Mult_Buf[65].Feature_n = FeatureBuf_163;
         Mult_Buf[65].Weight_n = Wgt_5_163;
         Mult_Buf[66].Feature_n = FeatureBuf_164;
         Mult_Buf[66].Weight_n = Wgt_5_164;
         Mult_Buf[67].Feature_n = FeatureBuf_165;
         Mult_Buf[67].Weight_n = Wgt_5_165;
         Mult_Buf[68].Feature_n = FeatureBuf_166;
         Mult_Buf[68].Weight_n = Wgt_5_166;
         Mult_Buf[69].Feature_n = FeatureBuf_167;
         Mult_Buf[69].Weight_n = Wgt_5_167;
         Mult_Buf[70].Feature_n = FeatureBuf_168;
         Mult_Buf[70].Weight_n = Wgt_5_168;
         Mult_Buf[71].Feature_n = FeatureBuf_169;
         Mult_Buf[71].Weight_n = Wgt_5_169;
         Mult_Buf[72].Feature_n = FeatureBuf_170;
         Mult_Buf[72].Weight_n = Wgt_5_170;
         Mult_Buf[73].Feature_n = FeatureBuf_171;
         Mult_Buf[73].Weight_n = Wgt_5_171;
         Mult_Buf[74].Feature_n = FeatureBuf_172;
         Mult_Buf[74].Weight_n = Wgt_5_172;
         Mult_Buf[75].Feature_n = FeatureBuf_173;
         Mult_Buf[75].Weight_n = Wgt_5_173;
         Mult_Buf[76].Feature_n = FeatureBuf_174;
         Mult_Buf[76].Weight_n = Wgt_5_174;
         Mult_Buf[77].Feature_n = FeatureBuf_175;
         Mult_Buf[77].Weight_n = Wgt_5_175;
         Mult_Buf[78].Feature_n = FeatureBuf_176;
         Mult_Buf[78].Weight_n = Wgt_5_176;
         Mult_Buf[79].Feature_n = FeatureBuf_177;
         Mult_Buf[79].Weight_n = Wgt_5_177;
         Mult_Buf[80].Feature_n = FeatureBuf_178;
         Mult_Buf[80].Weight_n = Wgt_5_178;
         Mult_Buf[81].Feature_n = FeatureBuf_179;
         Mult_Buf[81].Weight_n = Wgt_5_179;
         Mult_Buf[82].Feature_n = FeatureBuf_180;
         Mult_Buf[82].Weight_n = Wgt_5_180;
         Mult_Buf[83].Feature_n = FeatureBuf_181;
         Mult_Buf[83].Weight_n = Wgt_5_181;
         Mult_Buf[84].Feature_n = FeatureBuf_182;
         Mult_Buf[84].Weight_n = Wgt_5_182;
         Mult_Buf[85].Feature_n = FeatureBuf_183;
         Mult_Buf[85].Weight_n = Wgt_5_183;
         Mult_Buf[86].Feature_n = FeatureBuf_184;
         Mult_Buf[86].Weight_n = Wgt_5_184;
         Mult_Buf[87].Feature_n = FeatureBuf_185;
         Mult_Buf[87].Weight_n = Wgt_5_185;
         Mult_Buf[88].Feature_n = FeatureBuf_186;
         Mult_Buf[88].Weight_n = Wgt_5_186;
         Mult_Buf[89].Feature_n = FeatureBuf_187;
         Mult_Buf[89].Weight_n = Wgt_5_187;
         Mult_Buf[90].Feature_n = FeatureBuf_188;
         Mult_Buf[90].Weight_n = Wgt_5_188;
         Mult_Buf[91].Feature_n = FeatureBuf_189;
         Mult_Buf[91].Weight_n = Wgt_5_189;
         Mult_Buf[92].Feature_n = FeatureBuf_190;
         Mult_Buf[92].Weight_n = Wgt_5_190;
         Mult_Buf[93].Feature_n = FeatureBuf_191;
         Mult_Buf[93].Weight_n = Wgt_5_191;
         Mult_Buf[94].Feature_n = FeatureBuf_192;
         Mult_Buf[94].Weight_n = Wgt_5_192;
         Mult_Buf[95].Feature_n = FeatureBuf_193;
         Mult_Buf[95].Weight_n = Wgt_5_193;
         Mult_Buf[96].Feature_n = FeatureBuf_194;
         Mult_Buf[96].Weight_n = Wgt_5_194;
         Mult_Buf[97].Feature_n = FeatureBuf_195;
         Mult_Buf[97].Weight_n = Wgt_5_195;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     //Collect Partial result form Adder
         Res_2_3_n = Part_Res;
     end
    44:begin
     nxt_state = 45;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_196;
         Mult_Buf[0].Weight_n = Wgt_5_196;
         Mult_Buf[1].Feature_n = FeatureBuf_197;
         Mult_Buf[1].Weight_n = Wgt_5_197;
         Mult_Buf[2].Feature_n = FeatureBuf_198;
         Mult_Buf[2].Weight_n = Wgt_5_198;
         Mult_Buf[3].Feature_n = FeatureBuf_199;
         Mult_Buf[3].Weight_n = Wgt_5_199;
         Mult_Buf[4].Feature_n = FeatureBuf_200;
         Mult_Buf[4].Weight_n = Wgt_5_200;
         Mult_Buf[5].Feature_n = FeatureBuf_201;
         Mult_Buf[5].Weight_n = Wgt_5_201;
         Mult_Buf[6].Feature_n = FeatureBuf_202;
         Mult_Buf[6].Weight_n = Wgt_5_202;
         Mult_Buf[7].Feature_n = FeatureBuf_203;
         Mult_Buf[7].Weight_n = Wgt_5_203;
         Mult_Buf[8].Feature_n = FeatureBuf_204;
         Mult_Buf[8].Weight_n = Wgt_5_204;
         Mult_Buf[9].Feature_n = FeatureBuf_205;
         Mult_Buf[9].Weight_n = Wgt_5_205;
         Mult_Buf[10].Feature_n = FeatureBuf_206;
         Mult_Buf[10].Weight_n = Wgt_5_206;
         Mult_Buf[11].Feature_n = FeatureBuf_207;
         Mult_Buf[11].Weight_n = Wgt_5_207;
         Mult_Buf[12].Feature_n = FeatureBuf_208;
         Mult_Buf[12].Weight_n = Wgt_5_208;
         Mult_Buf[13].Feature_n = FeatureBuf_209;
         Mult_Buf[13].Weight_n = Wgt_5_209;
         Mult_Buf[14].Feature_n = FeatureBuf_210;
         Mult_Buf[14].Weight_n = Wgt_5_210;
         Mult_Buf[15].Feature_n = FeatureBuf_211;
         Mult_Buf[15].Weight_n = Wgt_5_211;
         Mult_Buf[16].Feature_n = FeatureBuf_212;
         Mult_Buf[16].Weight_n = Wgt_5_212;
         Mult_Buf[17].Feature_n = FeatureBuf_213;
         Mult_Buf[17].Weight_n = Wgt_5_213;
         Mult_Buf[18].Feature_n = FeatureBuf_214;
         Mult_Buf[18].Weight_n = Wgt_5_214;
         Mult_Buf[19].Feature_n = FeatureBuf_215;
         Mult_Buf[19].Weight_n = Wgt_5_215;
         Mult_Buf[20].Feature_n = FeatureBuf_216;
         Mult_Buf[20].Weight_n = Wgt_5_216;
         Mult_Buf[21].Feature_n = FeatureBuf_217;
         Mult_Buf[21].Weight_n = Wgt_5_217;
         Mult_Buf[22].Feature_n = FeatureBuf_218;
         Mult_Buf[22].Weight_n = Wgt_5_218;
         Mult_Buf[23].Feature_n = FeatureBuf_219;
         Mult_Buf[23].Weight_n = Wgt_5_219;
         Mult_Buf[24].Feature_n = FeatureBuf_220;
         Mult_Buf[24].Weight_n = Wgt_5_220;
         Mult_Buf[25].Feature_n = FeatureBuf_221;
         Mult_Buf[25].Weight_n = Wgt_5_221;
         Mult_Buf[26].Feature_n = FeatureBuf_222;
         Mult_Buf[26].Weight_n = Wgt_5_222;
         Mult_Buf[27].Feature_n = FeatureBuf_223;
         Mult_Buf[27].Weight_n = Wgt_5_223;
         Mult_Buf[28].Feature_n = FeatureBuf_224;
         Mult_Buf[28].Weight_n = Wgt_5_224;
         Mult_Buf[29].Feature_n = FeatureBuf_225;
         Mult_Buf[29].Weight_n = Wgt_5_225;
         Mult_Buf[30].Feature_n = FeatureBuf_226;
         Mult_Buf[30].Weight_n = Wgt_5_226;
         Mult_Buf[31].Feature_n = FeatureBuf_227;
         Mult_Buf[31].Weight_n = Wgt_5_227;
         Mult_Buf[32].Feature_n = FeatureBuf_228;
         Mult_Buf[32].Weight_n = Wgt_5_228;
         Mult_Buf[33].Feature_n = FeatureBuf_229;
         Mult_Buf[33].Weight_n = Wgt_5_229;
         Mult_Buf[34].Feature_n = FeatureBuf_230;
         Mult_Buf[34].Weight_n = Wgt_5_230;
         Mult_Buf[35].Feature_n = FeatureBuf_231;
         Mult_Buf[35].Weight_n = Wgt_5_231;
         Mult_Buf[36].Feature_n = FeatureBuf_232;
         Mult_Buf[36].Weight_n = Wgt_5_232;
         Mult_Buf[37].Feature_n = FeatureBuf_233;
         Mult_Buf[37].Weight_n = Wgt_5_233;
         Mult_Buf[38].Feature_n = FeatureBuf_234;
         Mult_Buf[38].Weight_n = Wgt_5_234;
         Mult_Buf[39].Feature_n = FeatureBuf_235;
         Mult_Buf[39].Weight_n = Wgt_5_235;
         Mult_Buf[40].Feature_n = FeatureBuf_236;
         Mult_Buf[40].Weight_n = Wgt_5_236;
         Mult_Buf[41].Feature_n = FeatureBuf_237;
         Mult_Buf[41].Weight_n = Wgt_5_237;
         Mult_Buf[42].Feature_n = FeatureBuf_238;
         Mult_Buf[42].Weight_n = Wgt_5_238;
         Mult_Buf[43].Feature_n = FeatureBuf_239;
         Mult_Buf[43].Weight_n = Wgt_5_239;
         Mult_Buf[44].Feature_n = FeatureBuf_240;
         Mult_Buf[44].Weight_n = Wgt_5_240;
         Mult_Buf[45].Feature_n = FeatureBuf_241;
         Mult_Buf[45].Weight_n = Wgt_5_241;
         Mult_Buf[46].Feature_n = FeatureBuf_242;
         Mult_Buf[46].Weight_n = Wgt_5_242;
         Mult_Buf[47].Feature_n = FeatureBuf_243;
         Mult_Buf[47].Weight_n = Wgt_5_243;
         Mult_Buf[48].Feature_n = FeatureBuf_244;
         Mult_Buf[48].Weight_n = Wgt_5_244;
         Mult_Buf[49].Feature_n = FeatureBuf_245;
         Mult_Buf[49].Weight_n = Wgt_5_245;
         Mult_Buf[50].Feature_n = FeatureBuf_246;
         Mult_Buf[50].Weight_n = Wgt_5_246;
         Mult_Buf[51].Feature_n = FeatureBuf_247;
         Mult_Buf[51].Weight_n = Wgt_5_247;
         Mult_Buf[52].Feature_n = FeatureBuf_248;
         Mult_Buf[52].Weight_n = Wgt_5_248;
         Mult_Buf[53].Feature_n = FeatureBuf_249;
         Mult_Buf[53].Weight_n = Wgt_5_249;
         Mult_Buf[54].Feature_n = FeatureBuf_250;
         Mult_Buf[54].Weight_n = Wgt_5_250;
         Mult_Buf[55].Feature_n = FeatureBuf_251;
         Mult_Buf[55].Weight_n = Wgt_5_251;
         Mult_Buf[56].Feature_n = FeatureBuf_252;
         Mult_Buf[56].Weight_n = Wgt_5_252;
         Mult_Buf[57].Feature_n = FeatureBuf_253;
         Mult_Buf[57].Weight_n = Wgt_5_253;
         Mult_Buf[58].Feature_n = FeatureBuf_254;
         Mult_Buf[58].Weight_n = Wgt_5_254;
         Mult_Buf[59].Feature_n = FeatureBuf_255;
         Mult_Buf[59].Weight_n = Wgt_5_255;
         Mult_Buf[60].Feature_n = FeatureBuf_256;
         Mult_Buf[60].Weight_n = Wgt_5_256;
         Mult_Buf[61].Feature_n = FeatureBuf_257;
         Mult_Buf[61].Weight_n = Wgt_5_257;
         Mult_Buf[62].Feature_n = FeatureBuf_258;
         Mult_Buf[62].Weight_n = Wgt_5_258;
         Mult_Buf[63].Feature_n = FeatureBuf_259;
         Mult_Buf[63].Weight_n = Wgt_5_259;
         Mult_Buf[64].Feature_n = FeatureBuf_260;
         Mult_Buf[64].Weight_n = Wgt_5_260;
         Mult_Buf[65].Feature_n = FeatureBuf_261;
         Mult_Buf[65].Weight_n = Wgt_5_261;
         Mult_Buf[66].Feature_n = FeatureBuf_262;
         Mult_Buf[66].Weight_n = Wgt_5_262;
         Mult_Buf[67].Feature_n = FeatureBuf_263;
         Mult_Buf[67].Weight_n = Wgt_5_263;
         Mult_Buf[68].Feature_n = FeatureBuf_264;
         Mult_Buf[68].Weight_n = Wgt_5_264;
         Mult_Buf[69].Feature_n = FeatureBuf_265;
         Mult_Buf[69].Weight_n = Wgt_5_265;
         Mult_Buf[70].Feature_n = FeatureBuf_266;
         Mult_Buf[70].Weight_n = Wgt_5_266;
         Mult_Buf[71].Feature_n = FeatureBuf_267;
         Mult_Buf[71].Weight_n = Wgt_5_267;
         Mult_Buf[72].Feature_n = FeatureBuf_268;
         Mult_Buf[72].Weight_n = Wgt_5_268;
         Mult_Buf[73].Feature_n = FeatureBuf_269;
         Mult_Buf[73].Weight_n = Wgt_5_269;
         Mult_Buf[74].Feature_n = FeatureBuf_270;
         Mult_Buf[74].Weight_n = Wgt_5_270;
         Mult_Buf[75].Feature_n = FeatureBuf_271;
         Mult_Buf[75].Weight_n = Wgt_5_271;
         Mult_Buf[76].Feature_n = FeatureBuf_272;
         Mult_Buf[76].Weight_n = Wgt_5_272;
         Mult_Buf[77].Feature_n = FeatureBuf_273;
         Mult_Buf[77].Weight_n = Wgt_5_273;
         Mult_Buf[78].Feature_n = FeatureBuf_274;
         Mult_Buf[78].Weight_n = Wgt_5_274;
         Mult_Buf[79].Feature_n = FeatureBuf_275;
         Mult_Buf[79].Weight_n = Wgt_5_275;
         Mult_Buf[80].Feature_n = FeatureBuf_276;
         Mult_Buf[80].Weight_n = Wgt_5_276;
         Mult_Buf[81].Feature_n = FeatureBuf_277;
         Mult_Buf[81].Weight_n = Wgt_5_277;
         Mult_Buf[82].Feature_n = FeatureBuf_278;
         Mult_Buf[82].Weight_n = Wgt_5_278;
         Mult_Buf[83].Feature_n = FeatureBuf_279;
         Mult_Buf[83].Weight_n = Wgt_5_279;
         Mult_Buf[84].Feature_n = FeatureBuf_280;
         Mult_Buf[84].Weight_n = Wgt_5_280;
         Mult_Buf[85].Feature_n = FeatureBuf_281;
         Mult_Buf[85].Weight_n = Wgt_5_281;
         Mult_Buf[86].Feature_n = FeatureBuf_282;
         Mult_Buf[86].Weight_n = Wgt_5_282;
         Mult_Buf[87].Feature_n = FeatureBuf_283;
         Mult_Buf[87].Weight_n = Wgt_5_283;
         Mult_Buf[88].Feature_n = FeatureBuf_284;
         Mult_Buf[88].Weight_n = Wgt_5_284;
         Mult_Buf[89].Feature_n = FeatureBuf_285;
         Mult_Buf[89].Weight_n = Wgt_5_285;
         Mult_Buf[90].Feature_n = FeatureBuf_286;
         Mult_Buf[90].Weight_n = Wgt_5_286;
         Mult_Buf[91].Feature_n = FeatureBuf_287;
         Mult_Buf[91].Weight_n = Wgt_5_287;
         Mult_Buf[92].Feature_n = FeatureBuf_288;
         Mult_Buf[92].Weight_n = Wgt_5_288;
         Mult_Buf[93].Feature_n = FeatureBuf_289;
         Mult_Buf[93].Weight_n = Wgt_5_289;
         Mult_Buf[94].Feature_n = FeatureBuf_290;
         Mult_Buf[94].Weight_n = Wgt_5_290;
         Mult_Buf[95].Feature_n = FeatureBuf_291;
         Mult_Buf[95].Weight_n = Wgt_5_291;
         Mult_Buf[96].Feature_n = FeatureBuf_292;
         Mult_Buf[96].Weight_n = Wgt_5_292;
         Mult_Buf[97].Feature_n = FeatureBuf_293;
         Mult_Buf[97].Weight_n = Wgt_5_293;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     //Collect Partial result form Adder
         Res_2_4_n = Part_Res;
     end
    45:begin
     nxt_state = 46;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_294;
         Mult_Buf[0].Weight_n = Wgt_5_294;
         Mult_Buf[1].Feature_n = FeatureBuf_295;
         Mult_Buf[1].Weight_n = Wgt_5_295;
         Mult_Buf[2].Feature_n = FeatureBuf_296;
         Mult_Buf[2].Weight_n = Wgt_5_296;
         Mult_Buf[3].Feature_n = FeatureBuf_297;
         Mult_Buf[3].Weight_n = Wgt_5_297;
         Mult_Buf[4].Feature_n = FeatureBuf_298;
         Mult_Buf[4].Weight_n = Wgt_5_298;
         Mult_Buf[5].Feature_n = FeatureBuf_299;
         Mult_Buf[5].Weight_n = Wgt_5_299;
         Mult_Buf[6].Feature_n = FeatureBuf_300;
         Mult_Buf[6].Weight_n = Wgt_5_300;
         Mult_Buf[7].Feature_n = FeatureBuf_301;
         Mult_Buf[7].Weight_n = Wgt_5_301;
         Mult_Buf[8].Feature_n = FeatureBuf_302;
         Mult_Buf[8].Weight_n = Wgt_5_302;
         Mult_Buf[9].Feature_n = FeatureBuf_303;
         Mult_Buf[9].Weight_n = Wgt_5_303;
         Mult_Buf[10].Feature_n = FeatureBuf_304;
         Mult_Buf[10].Weight_n = Wgt_5_304;
         Mult_Buf[11].Feature_n = FeatureBuf_305;
         Mult_Buf[11].Weight_n = Wgt_5_305;
         Mult_Buf[12].Feature_n = FeatureBuf_306;
         Mult_Buf[12].Weight_n = Wgt_5_306;
         Mult_Buf[13].Feature_n = FeatureBuf_307;
         Mult_Buf[13].Weight_n = Wgt_5_307;
         Mult_Buf[14].Feature_n = FeatureBuf_308;
         Mult_Buf[14].Weight_n = Wgt_5_308;
         Mult_Buf[15].Feature_n = FeatureBuf_309;
         Mult_Buf[15].Weight_n = Wgt_5_309;
         Mult_Buf[16].Feature_n = FeatureBuf_310;
         Mult_Buf[16].Weight_n = Wgt_5_310;
         Mult_Buf[17].Feature_n = FeatureBuf_311;
         Mult_Buf[17].Weight_n = Wgt_5_311;
         Mult_Buf[18].Feature_n = FeatureBuf_312;
         Mult_Buf[18].Weight_n = Wgt_5_312;
         Mult_Buf[19].Feature_n = FeatureBuf_313;
         Mult_Buf[19].Weight_n = Wgt_5_313;
         Mult_Buf[20].Feature_n = FeatureBuf_314;
         Mult_Buf[20].Weight_n = Wgt_5_314;
         Mult_Buf[21].Feature_n = FeatureBuf_315;
         Mult_Buf[21].Weight_n = Wgt_5_315;
         Mult_Buf[22].Feature_n = FeatureBuf_316;
         Mult_Buf[22].Weight_n = Wgt_5_316;
         Mult_Buf[23].Feature_n = FeatureBuf_317;
         Mult_Buf[23].Weight_n = Wgt_5_317;
         Mult_Buf[24].Feature_n = FeatureBuf_318;
         Mult_Buf[24].Weight_n = Wgt_5_318;
         Mult_Buf[25].Feature_n = FeatureBuf_319;
         Mult_Buf[25].Weight_n = Wgt_5_319;
         Mult_Buf[26].Feature_n = FeatureBuf_320;
         Mult_Buf[26].Weight_n = Wgt_5_320;
         Mult_Buf[27].Feature_n = FeatureBuf_321;
         Mult_Buf[27].Weight_n = Wgt_5_321;
         Mult_Buf[28].Feature_n = FeatureBuf_322;
         Mult_Buf[28].Weight_n = Wgt_5_322;
         Mult_Buf[29].Feature_n = FeatureBuf_323;
         Mult_Buf[29].Weight_n = Wgt_5_323;
         Mult_Buf[30].Feature_n = FeatureBuf_324;
         Mult_Buf[30].Weight_n = Wgt_5_324;
         Mult_Buf[31].Feature_n = FeatureBuf_325;
         Mult_Buf[31].Weight_n = Wgt_5_325;
         Mult_Buf[32].Feature_n = FeatureBuf_326;
         Mult_Buf[32].Weight_n = Wgt_5_326;
         Mult_Buf[33].Feature_n = FeatureBuf_327;
         Mult_Buf[33].Weight_n = Wgt_5_327;
         Mult_Buf[34].Feature_n = FeatureBuf_328;
         Mult_Buf[34].Weight_n = Wgt_5_328;
         Mult_Buf[35].Feature_n = FeatureBuf_329;
         Mult_Buf[35].Weight_n = Wgt_5_329;
         Mult_Buf[36].Feature_n = FeatureBuf_330;
         Mult_Buf[36].Weight_n = Wgt_5_330;
         Mult_Buf[37].Feature_n = FeatureBuf_331;
         Mult_Buf[37].Weight_n = Wgt_5_331;
         Mult_Buf[38].Feature_n = FeatureBuf_332;
         Mult_Buf[38].Weight_n = Wgt_5_332;
         Mult_Buf[39].Feature_n = FeatureBuf_333;
         Mult_Buf[39].Weight_n = Wgt_5_333;
         Mult_Buf[40].Feature_n = FeatureBuf_334;
         Mult_Buf[40].Weight_n = Wgt_5_334;
         Mult_Buf[41].Feature_n = FeatureBuf_335;
         Mult_Buf[41].Weight_n = Wgt_5_335;
         Mult_Buf[42].Feature_n = FeatureBuf_336;
         Mult_Buf[42].Weight_n = Wgt_5_336;
         Mult_Buf[43].Feature_n = FeatureBuf_337;
         Mult_Buf[43].Weight_n = Wgt_5_337;
         Mult_Buf[44].Feature_n = FeatureBuf_338;
         Mult_Buf[44].Weight_n = Wgt_5_338;
         Mult_Buf[45].Feature_n = FeatureBuf_339;
         Mult_Buf[45].Weight_n = Wgt_5_339;
         Mult_Buf[46].Feature_n = FeatureBuf_340;
         Mult_Buf[46].Weight_n = Wgt_5_340;
         Mult_Buf[47].Feature_n = FeatureBuf_341;
         Mult_Buf[47].Weight_n = Wgt_5_341;
         Mult_Buf[48].Feature_n = FeatureBuf_342;
         Mult_Buf[48].Weight_n = Wgt_5_342;
         Mult_Buf[49].Feature_n = FeatureBuf_343;
         Mult_Buf[49].Weight_n = Wgt_5_343;
         Mult_Buf[50].Feature_n = FeatureBuf_344;
         Mult_Buf[50].Weight_n = Wgt_5_344;
         Mult_Buf[51].Feature_n = FeatureBuf_345;
         Mult_Buf[51].Weight_n = Wgt_5_345;
         Mult_Buf[52].Feature_n = FeatureBuf_346;
         Mult_Buf[52].Weight_n = Wgt_5_346;
         Mult_Buf[53].Feature_n = FeatureBuf_347;
         Mult_Buf[53].Weight_n = Wgt_5_347;
         Mult_Buf[54].Feature_n = FeatureBuf_348;
         Mult_Buf[54].Weight_n = Wgt_5_348;
         Mult_Buf[55].Feature_n = FeatureBuf_349;
         Mult_Buf[55].Weight_n = Wgt_5_349;
         Mult_Buf[56].Feature_n = FeatureBuf_350;
         Mult_Buf[56].Weight_n = Wgt_5_350;
         Mult_Buf[57].Feature_n = FeatureBuf_351;
         Mult_Buf[57].Weight_n = Wgt_5_351;
         Mult_Buf[58].Feature_n = FeatureBuf_352;
         Mult_Buf[58].Weight_n = Wgt_5_352;
         Mult_Buf[59].Feature_n = FeatureBuf_353;
         Mult_Buf[59].Weight_n = Wgt_5_353;
         Mult_Buf[60].Feature_n = FeatureBuf_354;
         Mult_Buf[60].Weight_n = Wgt_5_354;
         Mult_Buf[61].Feature_n = FeatureBuf_355;
         Mult_Buf[61].Weight_n = Wgt_5_355;
         Mult_Buf[62].Feature_n = FeatureBuf_356;
         Mult_Buf[62].Weight_n = Wgt_5_356;
         Mult_Buf[63].Feature_n = FeatureBuf_357;
         Mult_Buf[63].Weight_n = Wgt_5_357;
         Mult_Buf[64].Feature_n = FeatureBuf_358;
         Mult_Buf[64].Weight_n = Wgt_5_358;
         Mult_Buf[65].Feature_n = FeatureBuf_359;
         Mult_Buf[65].Weight_n = Wgt_5_359;
         Mult_Buf[66].Feature_n = FeatureBuf_360;
         Mult_Buf[66].Weight_n = Wgt_5_360;
         Mult_Buf[67].Feature_n = FeatureBuf_361;
         Mult_Buf[67].Weight_n = Wgt_5_361;
         Mult_Buf[68].Feature_n = FeatureBuf_362;
         Mult_Buf[68].Weight_n = Wgt_5_362;
         Mult_Buf[69].Feature_n = FeatureBuf_363;
         Mult_Buf[69].Weight_n = Wgt_5_363;
         Mult_Buf[70].Feature_n = FeatureBuf_364;
         Mult_Buf[70].Weight_n = Wgt_5_364;
         Mult_Buf[71].Feature_n = FeatureBuf_365;
         Mult_Buf[71].Weight_n = Wgt_5_365;
         Mult_Buf[72].Feature_n = FeatureBuf_366;
         Mult_Buf[72].Weight_n = Wgt_5_366;
         Mult_Buf[73].Feature_n = FeatureBuf_367;
         Mult_Buf[73].Weight_n = Wgt_5_367;
         Mult_Buf[74].Feature_n = FeatureBuf_368;
         Mult_Buf[74].Weight_n = Wgt_5_368;
         Mult_Buf[75].Feature_n = FeatureBuf_369;
         Mult_Buf[75].Weight_n = Wgt_5_369;
         Mult_Buf[76].Feature_n = FeatureBuf_370;
         Mult_Buf[76].Weight_n = Wgt_5_370;
         Mult_Buf[77].Feature_n = FeatureBuf_371;
         Mult_Buf[77].Weight_n = Wgt_5_371;
         Mult_Buf[78].Feature_n = FeatureBuf_372;
         Mult_Buf[78].Weight_n = Wgt_5_372;
         Mult_Buf[79].Feature_n = FeatureBuf_373;
         Mult_Buf[79].Weight_n = Wgt_5_373;
         Mult_Buf[80].Feature_n = FeatureBuf_374;
         Mult_Buf[80].Weight_n = Wgt_5_374;
         Mult_Buf[81].Feature_n = FeatureBuf_375;
         Mult_Buf[81].Weight_n = Wgt_5_375;
         Mult_Buf[82].Feature_n = FeatureBuf_376;
         Mult_Buf[82].Weight_n = Wgt_5_376;
         Mult_Buf[83].Feature_n = FeatureBuf_377;
         Mult_Buf[83].Weight_n = Wgt_5_377;
         Mult_Buf[84].Feature_n = FeatureBuf_378;
         Mult_Buf[84].Weight_n = Wgt_5_378;
         Mult_Buf[85].Feature_n = FeatureBuf_379;
         Mult_Buf[85].Weight_n = Wgt_5_379;
         Mult_Buf[86].Feature_n = FeatureBuf_380;
         Mult_Buf[86].Weight_n = Wgt_5_380;
         Mult_Buf[87].Feature_n = FeatureBuf_381;
         Mult_Buf[87].Weight_n = Wgt_5_381;
         Mult_Buf[88].Feature_n = FeatureBuf_382;
         Mult_Buf[88].Weight_n = Wgt_5_382;
         Mult_Buf[89].Feature_n = FeatureBuf_383;
         Mult_Buf[89].Weight_n = Wgt_5_383;
         Mult_Buf[90].Feature_n = FeatureBuf_384;
         Mult_Buf[90].Weight_n = Wgt_5_384;
         Mult_Buf[91].Feature_n = FeatureBuf_385;
         Mult_Buf[91].Weight_n = Wgt_5_385;
         Mult_Buf[92].Feature_n = FeatureBuf_386;
         Mult_Buf[92].Weight_n = Wgt_5_386;
         Mult_Buf[93].Feature_n = FeatureBuf_387;
         Mult_Buf[93].Weight_n = Wgt_5_387;
         Mult_Buf[94].Feature_n = FeatureBuf_388;
         Mult_Buf[94].Weight_n = Wgt_5_388;
         Mult_Buf[95].Feature_n = FeatureBuf_389;
         Mult_Buf[95].Weight_n = Wgt_5_389;
         Mult_Buf[96].Feature_n = FeatureBuf_390;
         Mult_Buf[96].Weight_n = Wgt_5_390;
         Mult_Buf[97].Feature_n = FeatureBuf_391;
         Mult_Buf[97].Weight_n = Wgt_5_391;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     //Collect Partial result form Adder
         Res_2_5_n = Part_Res;
     //Collect result from final Adder
         Res1_n = Final_Res;
     end
    46:begin
     nxt_state = 47;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_392;
         Mult_Buf[0].Weight_n = Wgt_5_392;
         Mult_Buf[1].Feature_n = FeatureBuf_393;
         Mult_Buf[1].Weight_n = Wgt_5_393;
         Mult_Buf[2].Feature_n = FeatureBuf_394;
         Mult_Buf[2].Weight_n = Wgt_5_394;
         Mult_Buf[3].Feature_n = FeatureBuf_395;
         Mult_Buf[3].Weight_n = Wgt_5_395;
         Mult_Buf[4].Feature_n = FeatureBuf_396;
         Mult_Buf[4].Weight_n = Wgt_5_396;
         Mult_Buf[5].Feature_n = FeatureBuf_397;
         Mult_Buf[5].Weight_n = Wgt_5_397;
         Mult_Buf[6].Feature_n = FeatureBuf_398;
         Mult_Buf[6].Weight_n = Wgt_5_398;
         Mult_Buf[7].Feature_n = FeatureBuf_399;
         Mult_Buf[7].Weight_n = Wgt_5_399;
         Mult_Buf[8].Feature_n = FeatureBuf_400;
         Mult_Buf[8].Weight_n = Wgt_5_400;
         Mult_Buf[9].Feature_n = FeatureBuf_401;
         Mult_Buf[9].Weight_n = Wgt_5_401;
         Mult_Buf[10].Feature_n = FeatureBuf_402;
         Mult_Buf[10].Weight_n = Wgt_5_402;
         Mult_Buf[11].Feature_n = FeatureBuf_403;
         Mult_Buf[11].Weight_n = Wgt_5_403;
         Mult_Buf[12].Feature_n = FeatureBuf_404;
         Mult_Buf[12].Weight_n = Wgt_5_404;
         Mult_Buf[13].Feature_n = FeatureBuf_405;
         Mult_Buf[13].Weight_n = Wgt_5_405;
         Mult_Buf[14].Feature_n = FeatureBuf_406;
         Mult_Buf[14].Weight_n = Wgt_5_406;
         Mult_Buf[15].Feature_n = FeatureBuf_407;
         Mult_Buf[15].Weight_n = Wgt_5_407;
         Mult_Buf[16].Feature_n = FeatureBuf_408;
         Mult_Buf[16].Weight_n = Wgt_5_408;
         Mult_Buf[17].Feature_n = FeatureBuf_409;
         Mult_Buf[17].Weight_n = Wgt_5_409;
         Mult_Buf[18].Feature_n = FeatureBuf_410;
         Mult_Buf[18].Weight_n = Wgt_5_410;
         Mult_Buf[19].Feature_n = FeatureBuf_411;
         Mult_Buf[19].Weight_n = Wgt_5_411;
         Mult_Buf[20].Feature_n = FeatureBuf_412;
         Mult_Buf[20].Weight_n = Wgt_5_412;
         Mult_Buf[21].Feature_n = FeatureBuf_413;
         Mult_Buf[21].Weight_n = Wgt_5_413;
         Mult_Buf[22].Feature_n = FeatureBuf_414;
         Mult_Buf[22].Weight_n = Wgt_5_414;
         Mult_Buf[23].Feature_n = FeatureBuf_415;
         Mult_Buf[23].Weight_n = Wgt_5_415;
         Mult_Buf[24].Feature_n = FeatureBuf_416;
         Mult_Buf[24].Weight_n = Wgt_5_416;
         Mult_Buf[25].Feature_n = FeatureBuf_417;
         Mult_Buf[25].Weight_n = Wgt_5_417;
         Mult_Buf[26].Feature_n = FeatureBuf_418;
         Mult_Buf[26].Weight_n = Wgt_5_418;
         Mult_Buf[27].Feature_n = FeatureBuf_419;
         Mult_Buf[27].Weight_n = Wgt_5_419;
         Mult_Buf[28].Feature_n = FeatureBuf_420;
         Mult_Buf[28].Weight_n = Wgt_5_420;
         Mult_Buf[29].Feature_n = FeatureBuf_421;
         Mult_Buf[29].Weight_n = Wgt_5_421;
         Mult_Buf[30].Feature_n = FeatureBuf_422;
         Mult_Buf[30].Weight_n = Wgt_5_422;
         Mult_Buf[31].Feature_n = FeatureBuf_423;
         Mult_Buf[31].Weight_n = Wgt_5_423;
         Mult_Buf[32].Feature_n = FeatureBuf_424;
         Mult_Buf[32].Weight_n = Wgt_5_424;
         Mult_Buf[33].Feature_n = FeatureBuf_425;
         Mult_Buf[33].Weight_n = Wgt_5_425;
         Mult_Buf[34].Feature_n = FeatureBuf_426;
         Mult_Buf[34].Weight_n = Wgt_5_426;
         Mult_Buf[35].Feature_n = FeatureBuf_427;
         Mult_Buf[35].Weight_n = Wgt_5_427;
         Mult_Buf[36].Feature_n = FeatureBuf_428;
         Mult_Buf[36].Weight_n = Wgt_5_428;
         Mult_Buf[37].Feature_n = FeatureBuf_429;
         Mult_Buf[37].Weight_n = Wgt_5_429;
         Mult_Buf[38].Feature_n = FeatureBuf_430;
         Mult_Buf[38].Weight_n = Wgt_5_430;
         Mult_Buf[39].Feature_n = FeatureBuf_431;
         Mult_Buf[39].Weight_n = Wgt_5_431;
         Mult_Buf[40].Feature_n = FeatureBuf_432;
         Mult_Buf[40].Weight_n = Wgt_5_432;
         Mult_Buf[41].Feature_n = FeatureBuf_433;
         Mult_Buf[41].Weight_n = Wgt_5_433;
         Mult_Buf[42].Feature_n = FeatureBuf_434;
         Mult_Buf[42].Weight_n = Wgt_5_434;
         Mult_Buf[43].Feature_n = FeatureBuf_435;
         Mult_Buf[43].Weight_n = Wgt_5_435;
         Mult_Buf[44].Feature_n = FeatureBuf_436;
         Mult_Buf[44].Weight_n = Wgt_5_436;
         Mult_Buf[45].Feature_n = FeatureBuf_437;
         Mult_Buf[45].Weight_n = Wgt_5_437;
         Mult_Buf[46].Feature_n = FeatureBuf_438;
         Mult_Buf[46].Weight_n = Wgt_5_438;
         Mult_Buf[47].Feature_n = FeatureBuf_439;
         Mult_Buf[47].Weight_n = Wgt_5_439;
         Mult_Buf[48].Feature_n = FeatureBuf_440;
         Mult_Buf[48].Weight_n = Wgt_5_440;
         Mult_Buf[49].Feature_n = FeatureBuf_441;
         Mult_Buf[49].Weight_n = Wgt_5_441;
         Mult_Buf[50].Feature_n = FeatureBuf_442;
         Mult_Buf[50].Weight_n = Wgt_5_442;
         Mult_Buf[51].Feature_n = FeatureBuf_443;
         Mult_Buf[51].Weight_n = Wgt_5_443;
         Mult_Buf[52].Feature_n = FeatureBuf_444;
         Mult_Buf[52].Weight_n = Wgt_5_444;
         Mult_Buf[53].Feature_n = FeatureBuf_445;
         Mult_Buf[53].Weight_n = Wgt_5_445;
         Mult_Buf[54].Feature_n = FeatureBuf_446;
         Mult_Buf[54].Weight_n = Wgt_5_446;
         Mult_Buf[55].Feature_n = FeatureBuf_447;
         Mult_Buf[55].Weight_n = Wgt_5_447;
         Mult_Buf[56].Feature_n = FeatureBuf_448;
         Mult_Buf[56].Weight_n = Wgt_5_448;
         Mult_Buf[57].Feature_n = FeatureBuf_449;
         Mult_Buf[57].Weight_n = Wgt_5_449;
         Mult_Buf[58].Feature_n = FeatureBuf_450;
         Mult_Buf[58].Weight_n = Wgt_5_450;
         Mult_Buf[59].Feature_n = FeatureBuf_451;
         Mult_Buf[59].Weight_n = Wgt_5_451;
         Mult_Buf[60].Feature_n = FeatureBuf_452;
         Mult_Buf[60].Weight_n = Wgt_5_452;
         Mult_Buf[61].Feature_n = FeatureBuf_453;
         Mult_Buf[61].Weight_n = Wgt_5_453;
         Mult_Buf[62].Feature_n = FeatureBuf_454;
         Mult_Buf[62].Weight_n = Wgt_5_454;
         Mult_Buf[63].Feature_n = FeatureBuf_455;
         Mult_Buf[63].Weight_n = Wgt_5_455;
         Mult_Buf[64].Feature_n = FeatureBuf_456;
         Mult_Buf[64].Weight_n = Wgt_5_456;
         Mult_Buf[65].Feature_n = FeatureBuf_457;
         Mult_Buf[65].Weight_n = Wgt_5_457;
         Mult_Buf[66].Feature_n = FeatureBuf_458;
         Mult_Buf[66].Weight_n = Wgt_5_458;
         Mult_Buf[67].Feature_n = FeatureBuf_459;
         Mult_Buf[67].Weight_n = Wgt_5_459;
         Mult_Buf[68].Feature_n = FeatureBuf_460;
         Mult_Buf[68].Weight_n = Wgt_5_460;
         Mult_Buf[69].Feature_n = FeatureBuf_461;
         Mult_Buf[69].Weight_n = Wgt_5_461;
         Mult_Buf[70].Feature_n = FeatureBuf_462;
         Mult_Buf[70].Weight_n = Wgt_5_462;
         Mult_Buf[71].Feature_n = FeatureBuf_463;
         Mult_Buf[71].Weight_n = Wgt_5_463;
         Mult_Buf[72].Feature_n = FeatureBuf_464;
         Mult_Buf[72].Weight_n = Wgt_5_464;
         Mult_Buf[73].Feature_n = FeatureBuf_465;
         Mult_Buf[73].Weight_n = Wgt_5_465;
         Mult_Buf[74].Feature_n = FeatureBuf_466;
         Mult_Buf[74].Weight_n = Wgt_5_466;
         Mult_Buf[75].Feature_n = FeatureBuf_467;
         Mult_Buf[75].Weight_n = Wgt_5_467;
         Mult_Buf[76].Feature_n = FeatureBuf_468;
         Mult_Buf[76].Weight_n = Wgt_5_468;
         Mult_Buf[77].Feature_n = FeatureBuf_469;
         Mult_Buf[77].Weight_n = Wgt_5_469;
         Mult_Buf[78].Feature_n = FeatureBuf_470;
         Mult_Buf[78].Weight_n = Wgt_5_470;
         Mult_Buf[79].Feature_n = FeatureBuf_471;
         Mult_Buf[79].Weight_n = Wgt_5_471;
         Mult_Buf[80].Feature_n = FeatureBuf_472;
         Mult_Buf[80].Weight_n = Wgt_5_472;
         Mult_Buf[81].Feature_n = FeatureBuf_473;
         Mult_Buf[81].Weight_n = Wgt_5_473;
         Mult_Buf[82].Feature_n = FeatureBuf_474;
         Mult_Buf[82].Weight_n = Wgt_5_474;
         Mult_Buf[83].Feature_n = FeatureBuf_475;
         Mult_Buf[83].Weight_n = Wgt_5_475;
         Mult_Buf[84].Feature_n = FeatureBuf_476;
         Mult_Buf[84].Weight_n = Wgt_5_476;
         Mult_Buf[85].Feature_n = FeatureBuf_477;
         Mult_Buf[85].Weight_n = Wgt_5_477;
         Mult_Buf[86].Feature_n = FeatureBuf_478;
         Mult_Buf[86].Weight_n = Wgt_5_478;
         Mult_Buf[87].Feature_n = FeatureBuf_479;
         Mult_Buf[87].Weight_n = Wgt_5_479;
         Mult_Buf[88].Feature_n = FeatureBuf_480;
         Mult_Buf[88].Weight_n = Wgt_5_480;
         Mult_Buf[89].Feature_n = FeatureBuf_481;
         Mult_Buf[89].Weight_n = Wgt_5_481;
         Mult_Buf[90].Feature_n = FeatureBuf_482;
         Mult_Buf[90].Weight_n = Wgt_5_482;
         Mult_Buf[91].Feature_n = FeatureBuf_483;
         Mult_Buf[91].Weight_n = Wgt_5_483;
         Mult_Buf[92].Feature_n = FeatureBuf_484;
         Mult_Buf[92].Weight_n = Wgt_5_484;
         Mult_Buf[93].Feature_n = FeatureBuf_485;
         Mult_Buf[93].Weight_n = Wgt_5_485;
         Mult_Buf[94].Feature_n = FeatureBuf_486;
         Mult_Buf[94].Weight_n = Wgt_5_486;
         Mult_Buf[95].Feature_n = FeatureBuf_487;
         Mult_Buf[95].Weight_n = Wgt_5_487;
         Mult_Buf[96].Feature_n = FeatureBuf_488;
         Mult_Buf[96].Weight_n = Wgt_5_488;
         Mult_Buf[97].Feature_n = FeatureBuf_489;
         Mult_Buf[97].Weight_n = Wgt_5_489;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     //Collect Partial result form Adder
         Res_2_6_n = Part_Res;
     end
    47:begin
     nxt_state = 48;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_490;
         Mult_Buf[0].Weight_n = Wgt_5_490;
         Mult_Buf[1].Feature_n = FeatureBuf_491;
         Mult_Buf[1].Weight_n = Wgt_5_491;
         Mult_Buf[2].Feature_n = FeatureBuf_492;
         Mult_Buf[2].Weight_n = Wgt_5_492;
         Mult_Buf[3].Feature_n = FeatureBuf_493;
         Mult_Buf[3].Weight_n = Wgt_5_493;
         Mult_Buf[4].Feature_n = FeatureBuf_494;
         Mult_Buf[4].Weight_n = Wgt_5_494;
         Mult_Buf[5].Feature_n = FeatureBuf_495;
         Mult_Buf[5].Weight_n = Wgt_5_495;
         Mult_Buf[6].Feature_n = FeatureBuf_496;
         Mult_Buf[6].Weight_n = Wgt_5_496;
         Mult_Buf[7].Feature_n = FeatureBuf_497;
         Mult_Buf[7].Weight_n = Wgt_5_497;
         Mult_Buf[8].Feature_n = FeatureBuf_498;
         Mult_Buf[8].Weight_n = Wgt_5_498;
         Mult_Buf[9].Feature_n = FeatureBuf_499;
         Mult_Buf[9].Weight_n = Wgt_5_499;
         Mult_Buf[10].Feature_n = FeatureBuf_500;
         Mult_Buf[10].Weight_n = Wgt_5_500;
         Mult_Buf[11].Feature_n = FeatureBuf_501;
         Mult_Buf[11].Weight_n = Wgt_5_501;
         Mult_Buf[12].Feature_n = FeatureBuf_502;
         Mult_Buf[12].Weight_n = Wgt_5_502;
         Mult_Buf[13].Feature_n = FeatureBuf_503;
         Mult_Buf[13].Weight_n = Wgt_5_503;
         Mult_Buf[14].Feature_n = FeatureBuf_504;
         Mult_Buf[14].Weight_n = Wgt_5_504;
         Mult_Buf[15].Feature_n = FeatureBuf_505;
         Mult_Buf[15].Weight_n = Wgt_5_505;
         Mult_Buf[16].Feature_n = FeatureBuf_506;
         Mult_Buf[16].Weight_n = Wgt_5_506;
         Mult_Buf[17].Feature_n = FeatureBuf_507;
         Mult_Buf[17].Weight_n = Wgt_5_507;
         Mult_Buf[18].Feature_n = FeatureBuf_508;
         Mult_Buf[18].Weight_n = Wgt_5_508;
         Mult_Buf[19].Feature_n = FeatureBuf_509;
         Mult_Buf[19].Weight_n = Wgt_5_509;
         Mult_Buf[20].Feature_n = FeatureBuf_510;
         Mult_Buf[20].Weight_n = Wgt_5_510;
         Mult_Buf[21].Feature_n = FeatureBuf_511;
         Mult_Buf[21].Weight_n = Wgt_5_511;
         Mult_Buf[22].Feature_n = FeatureBuf_512;
         Mult_Buf[22].Weight_n = Wgt_5_512;
         Mult_Buf[23].Feature_n = FeatureBuf_513;
         Mult_Buf[23].Weight_n = Wgt_5_513;
         Mult_Buf[24].Feature_n = FeatureBuf_514;
         Mult_Buf[24].Weight_n = Wgt_5_514;
         Mult_Buf[25].Feature_n = FeatureBuf_515;
         Mult_Buf[25].Weight_n = Wgt_5_515;
         Mult_Buf[26].Feature_n = FeatureBuf_516;
         Mult_Buf[26].Weight_n = Wgt_5_516;
         Mult_Buf[27].Feature_n = FeatureBuf_517;
         Mult_Buf[27].Weight_n = Wgt_5_517;
         Mult_Buf[28].Feature_n = FeatureBuf_518;
         Mult_Buf[28].Weight_n = Wgt_5_518;
         Mult_Buf[29].Feature_n = FeatureBuf_519;
         Mult_Buf[29].Weight_n = Wgt_5_519;
         Mult_Buf[30].Feature_n = FeatureBuf_520;
         Mult_Buf[30].Weight_n = Wgt_5_520;
         Mult_Buf[31].Feature_n = FeatureBuf_521;
         Mult_Buf[31].Weight_n = Wgt_5_521;
         Mult_Buf[32].Feature_n = FeatureBuf_522;
         Mult_Buf[32].Weight_n = Wgt_5_522;
         Mult_Buf[33].Feature_n = FeatureBuf_523;
         Mult_Buf[33].Weight_n = Wgt_5_523;
         Mult_Buf[34].Feature_n = FeatureBuf_524;
         Mult_Buf[34].Weight_n = Wgt_5_524;
         Mult_Buf[35].Feature_n = FeatureBuf_525;
         Mult_Buf[35].Weight_n = Wgt_5_525;
         Mult_Buf[36].Feature_n = FeatureBuf_526;
         Mult_Buf[36].Weight_n = Wgt_5_526;
         Mult_Buf[37].Feature_n = FeatureBuf_527;
         Mult_Buf[37].Weight_n = Wgt_5_527;
         Mult_Buf[38].Feature_n = FeatureBuf_528;
         Mult_Buf[38].Weight_n = Wgt_5_528;
         Mult_Buf[39].Feature_n = FeatureBuf_529;
         Mult_Buf[39].Weight_n = Wgt_5_529;
         Mult_Buf[40].Feature_n = FeatureBuf_530;
         Mult_Buf[40].Weight_n = Wgt_5_530;
         Mult_Buf[41].Feature_n = FeatureBuf_531;
         Mult_Buf[41].Weight_n = Wgt_5_531;
         Mult_Buf[42].Feature_n = FeatureBuf_532;
         Mult_Buf[42].Weight_n = Wgt_5_532;
         Mult_Buf[43].Feature_n = FeatureBuf_533;
         Mult_Buf[43].Weight_n = Wgt_5_533;
         Mult_Buf[44].Feature_n = FeatureBuf_534;
         Mult_Buf[44].Weight_n = Wgt_5_534;
         Mult_Buf[45].Feature_n = FeatureBuf_535;
         Mult_Buf[45].Weight_n = Wgt_5_535;
         Mult_Buf[46].Feature_n = FeatureBuf_536;
         Mult_Buf[46].Weight_n = Wgt_5_536;
         Mult_Buf[47].Feature_n = FeatureBuf_537;
         Mult_Buf[47].Weight_n = Wgt_5_537;
         Mult_Buf[48].Feature_n = FeatureBuf_538;
         Mult_Buf[48].Weight_n = Wgt_5_538;
         Mult_Buf[49].Feature_n = FeatureBuf_539;
         Mult_Buf[49].Weight_n = Wgt_5_539;
         Mult_Buf[50].Feature_n = FeatureBuf_540;
         Mult_Buf[50].Weight_n = Wgt_5_540;
         Mult_Buf[51].Feature_n = FeatureBuf_541;
         Mult_Buf[51].Weight_n = Wgt_5_541;
         Mult_Buf[52].Feature_n = FeatureBuf_542;
         Mult_Buf[52].Weight_n = Wgt_5_542;
         Mult_Buf[53].Feature_n = FeatureBuf_543;
         Mult_Buf[53].Weight_n = Wgt_5_543;
         Mult_Buf[54].Feature_n = FeatureBuf_544;
         Mult_Buf[54].Weight_n = Wgt_5_544;
         Mult_Buf[55].Feature_n = FeatureBuf_545;
         Mult_Buf[55].Weight_n = Wgt_5_545;
         Mult_Buf[56].Feature_n = FeatureBuf_546;
         Mult_Buf[56].Weight_n = Wgt_5_546;
         Mult_Buf[57].Feature_n = FeatureBuf_547;
         Mult_Buf[57].Weight_n = Wgt_5_547;
         Mult_Buf[58].Feature_n = FeatureBuf_548;
         Mult_Buf[58].Weight_n = Wgt_5_548;
         Mult_Buf[59].Feature_n = FeatureBuf_549;
         Mult_Buf[59].Weight_n = Wgt_5_549;
         Mult_Buf[60].Feature_n = FeatureBuf_550;
         Mult_Buf[60].Weight_n = Wgt_5_550;
         Mult_Buf[61].Feature_n = FeatureBuf_551;
         Mult_Buf[61].Weight_n = Wgt_5_551;
         Mult_Buf[62].Feature_n = FeatureBuf_552;
         Mult_Buf[62].Weight_n = Wgt_5_552;
         Mult_Buf[63].Feature_n = FeatureBuf_553;
         Mult_Buf[63].Weight_n = Wgt_5_553;
         Mult_Buf[64].Feature_n = FeatureBuf_554;
         Mult_Buf[64].Weight_n = Wgt_5_554;
         Mult_Buf[65].Feature_n = FeatureBuf_555;
         Mult_Buf[65].Weight_n = Wgt_5_555;
         Mult_Buf[66].Feature_n = FeatureBuf_556;
         Mult_Buf[66].Weight_n = Wgt_5_556;
         Mult_Buf[67].Feature_n = FeatureBuf_557;
         Mult_Buf[67].Weight_n = Wgt_5_557;
         Mult_Buf[68].Feature_n = FeatureBuf_558;
         Mult_Buf[68].Weight_n = Wgt_5_558;
         Mult_Buf[69].Feature_n = FeatureBuf_559;
         Mult_Buf[69].Weight_n = Wgt_5_559;
         Mult_Buf[70].Feature_n = FeatureBuf_560;
         Mult_Buf[70].Weight_n = Wgt_5_560;
         Mult_Buf[71].Feature_n = FeatureBuf_561;
         Mult_Buf[71].Weight_n = Wgt_5_561;
         Mult_Buf[72].Feature_n = FeatureBuf_562;
         Mult_Buf[72].Weight_n = Wgt_5_562;
         Mult_Buf[73].Feature_n = FeatureBuf_563;
         Mult_Buf[73].Weight_n = Wgt_5_563;
         Mult_Buf[74].Feature_n = FeatureBuf_564;
         Mult_Buf[74].Weight_n = Wgt_5_564;
         Mult_Buf[75].Feature_n = FeatureBuf_565;
         Mult_Buf[75].Weight_n = Wgt_5_565;
         Mult_Buf[76].Feature_n = FeatureBuf_566;
         Mult_Buf[76].Weight_n = Wgt_5_566;
         Mult_Buf[77].Feature_n = FeatureBuf_567;
         Mult_Buf[77].Weight_n = Wgt_5_567;
         Mult_Buf[78].Feature_n = FeatureBuf_568;
         Mult_Buf[78].Weight_n = Wgt_5_568;
         Mult_Buf[79].Feature_n = FeatureBuf_569;
         Mult_Buf[79].Weight_n = Wgt_5_569;
         Mult_Buf[80].Feature_n = FeatureBuf_570;
         Mult_Buf[80].Weight_n = Wgt_5_570;
         Mult_Buf[81].Feature_n = FeatureBuf_571;
         Mult_Buf[81].Weight_n = Wgt_5_571;
         Mult_Buf[82].Feature_n = FeatureBuf_572;
         Mult_Buf[82].Weight_n = Wgt_5_572;
         Mult_Buf[83].Feature_n = FeatureBuf_573;
         Mult_Buf[83].Weight_n = Wgt_5_573;
         Mult_Buf[84].Feature_n = FeatureBuf_574;
         Mult_Buf[84].Weight_n = Wgt_5_574;
         Mult_Buf[85].Feature_n = FeatureBuf_575;
         Mult_Buf[85].Weight_n = Wgt_5_575;
         Mult_Buf[86].Feature_n = FeatureBuf_576;
         Mult_Buf[86].Weight_n = Wgt_5_576;
         Mult_Buf[87].Feature_n = FeatureBuf_577;
         Mult_Buf[87].Weight_n = Wgt_5_577;
         Mult_Buf[88].Feature_n = FeatureBuf_578;
         Mult_Buf[88].Weight_n = Wgt_5_578;
         Mult_Buf[89].Feature_n = FeatureBuf_579;
         Mult_Buf[89].Weight_n = Wgt_5_579;
         Mult_Buf[90].Feature_n = FeatureBuf_580;
         Mult_Buf[90].Weight_n = Wgt_5_580;
         Mult_Buf[91].Feature_n = FeatureBuf_581;
         Mult_Buf[91].Weight_n = Wgt_5_581;
         Mult_Buf[92].Feature_n = FeatureBuf_582;
         Mult_Buf[92].Weight_n = Wgt_5_582;
         Mult_Buf[93].Feature_n = FeatureBuf_583;
         Mult_Buf[93].Weight_n = Wgt_5_583;
         Mult_Buf[94].Feature_n = FeatureBuf_584;
         Mult_Buf[94].Weight_n = Wgt_5_584;
         Mult_Buf[95].Feature_n = FeatureBuf_585;
         Mult_Buf[95].Weight_n = Wgt_5_585;
         Mult_Buf[96].Feature_n = FeatureBuf_586;
         Mult_Buf[96].Weight_n = Wgt_5_586;
         Mult_Buf[97].Feature_n = FeatureBuf_587;
         Mult_Buf[97].Weight_n = Wgt_5_587;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     //Collect Partial result form Adder
         Res_2_7_n = Part_Res;
     //Feed to final Adder
         A1 = Part_Res;
         A2 = Res_2_6_n;
         A3 = Res_2_5_n;
         A4 = Res_2_4_n;
         A5 = Res_2_3_n;
         A6 = Res_2_2_n;
         A7 = Res_2_1_n;
         A8 = Res_2_0_n;
     end
    48:begin
     nxt_state = 49;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_588;
         Mult_Buf[0].Weight_n = Wgt_5_588;
         Mult_Buf[1].Feature_n = FeatureBuf_589;
         Mult_Buf[1].Weight_n = Wgt_5_589;
         Mult_Buf[2].Feature_n = FeatureBuf_590;
         Mult_Buf[2].Weight_n = Wgt_5_590;
         Mult_Buf[3].Feature_n = FeatureBuf_591;
         Mult_Buf[3].Weight_n = Wgt_5_591;
         Mult_Buf[4].Feature_n = FeatureBuf_592;
         Mult_Buf[4].Weight_n = Wgt_5_592;
         Mult_Buf[5].Feature_n = FeatureBuf_593;
         Mult_Buf[5].Weight_n = Wgt_5_593;
         Mult_Buf[6].Feature_n = FeatureBuf_594;
         Mult_Buf[6].Weight_n = Wgt_5_594;
         Mult_Buf[7].Feature_n = FeatureBuf_595;
         Mult_Buf[7].Weight_n = Wgt_5_595;
         Mult_Buf[8].Feature_n = FeatureBuf_596;
         Mult_Buf[8].Weight_n = Wgt_5_596;
         Mult_Buf[9].Feature_n = FeatureBuf_597;
         Mult_Buf[9].Weight_n = Wgt_5_597;
         Mult_Buf[10].Feature_n = FeatureBuf_598;
         Mult_Buf[10].Weight_n = Wgt_5_598;
         Mult_Buf[11].Feature_n = FeatureBuf_599;
         Mult_Buf[11].Weight_n = Wgt_5_599;
         Mult_Buf[12].Feature_n = FeatureBuf_600;
         Mult_Buf[12].Weight_n = Wgt_5_600;
         Mult_Buf[13].Feature_n = FeatureBuf_601;
         Mult_Buf[13].Weight_n = Wgt_5_601;
         Mult_Buf[14].Feature_n = FeatureBuf_602;
         Mult_Buf[14].Weight_n = Wgt_5_602;
         Mult_Buf[15].Feature_n = FeatureBuf_603;
         Mult_Buf[15].Weight_n = Wgt_5_603;
         Mult_Buf[16].Feature_n = FeatureBuf_604;
         Mult_Buf[16].Weight_n = Wgt_5_604;
         Mult_Buf[17].Feature_n = FeatureBuf_605;
         Mult_Buf[17].Weight_n = Wgt_5_605;
         Mult_Buf[18].Feature_n = FeatureBuf_606;
         Mult_Buf[18].Weight_n = Wgt_5_606;
         Mult_Buf[19].Feature_n = FeatureBuf_607;
         Mult_Buf[19].Weight_n = Wgt_5_607;
         Mult_Buf[20].Feature_n = FeatureBuf_608;
         Mult_Buf[20].Weight_n = Wgt_5_608;
         Mult_Buf[21].Feature_n = FeatureBuf_609;
         Mult_Buf[21].Weight_n = Wgt_5_609;
         Mult_Buf[22].Feature_n = FeatureBuf_610;
         Mult_Buf[22].Weight_n = Wgt_5_610;
         Mult_Buf[23].Feature_n = FeatureBuf_611;
         Mult_Buf[23].Weight_n = Wgt_5_611;
         Mult_Buf[24].Feature_n = FeatureBuf_612;
         Mult_Buf[24].Weight_n = Wgt_5_612;
         Mult_Buf[25].Feature_n = FeatureBuf_613;
         Mult_Buf[25].Weight_n = Wgt_5_613;
         Mult_Buf[26].Feature_n = FeatureBuf_614;
         Mult_Buf[26].Weight_n = Wgt_5_614;
         Mult_Buf[27].Feature_n = FeatureBuf_615;
         Mult_Buf[27].Weight_n = Wgt_5_615;
         Mult_Buf[28].Feature_n = FeatureBuf_616;
         Mult_Buf[28].Weight_n = Wgt_5_616;
         Mult_Buf[29].Feature_n = FeatureBuf_617;
         Mult_Buf[29].Weight_n = Wgt_5_617;
         Mult_Buf[30].Feature_n = FeatureBuf_618;
         Mult_Buf[30].Weight_n = Wgt_5_618;
         Mult_Buf[31].Feature_n = FeatureBuf_619;
         Mult_Buf[31].Weight_n = Wgt_5_619;
         Mult_Buf[32].Feature_n = FeatureBuf_620;
         Mult_Buf[32].Weight_n = Wgt_5_620;
         Mult_Buf[33].Feature_n = FeatureBuf_621;
         Mult_Buf[33].Weight_n = Wgt_5_621;
         Mult_Buf[34].Feature_n = FeatureBuf_622;
         Mult_Buf[34].Weight_n = Wgt_5_622;
         Mult_Buf[35].Feature_n = FeatureBuf_623;
         Mult_Buf[35].Weight_n = Wgt_5_623;
         Mult_Buf[36].Feature_n = FeatureBuf_624;
         Mult_Buf[36].Weight_n = Wgt_5_624;
         Mult_Buf[37].Feature_n = FeatureBuf_625;
         Mult_Buf[37].Weight_n = Wgt_5_625;
         Mult_Buf[38].Feature_n = FeatureBuf_626;
         Mult_Buf[38].Weight_n = Wgt_5_626;
         Mult_Buf[39].Feature_n = FeatureBuf_627;
         Mult_Buf[39].Weight_n = Wgt_5_627;
         Mult_Buf[40].Feature_n = FeatureBuf_628;
         Mult_Buf[40].Weight_n = Wgt_5_628;
         Mult_Buf[41].Feature_n = FeatureBuf_629;
         Mult_Buf[41].Weight_n = Wgt_5_629;
         Mult_Buf[42].Feature_n = FeatureBuf_630;
         Mult_Buf[42].Weight_n = Wgt_5_630;
         Mult_Buf[43].Feature_n = FeatureBuf_631;
         Mult_Buf[43].Weight_n = Wgt_5_631;
         Mult_Buf[44].Feature_n = FeatureBuf_632;
         Mult_Buf[44].Weight_n = Wgt_5_632;
         Mult_Buf[45].Feature_n = FeatureBuf_633;
         Mult_Buf[45].Weight_n = Wgt_5_633;
         Mult_Buf[46].Feature_n = FeatureBuf_634;
         Mult_Buf[46].Weight_n = Wgt_5_634;
         Mult_Buf[47].Feature_n = FeatureBuf_635;
         Mult_Buf[47].Weight_n = Wgt_5_635;
         Mult_Buf[48].Feature_n = FeatureBuf_636;
         Mult_Buf[48].Weight_n = Wgt_5_636;
         Mult_Buf[49].Feature_n = FeatureBuf_637;
         Mult_Buf[49].Weight_n = Wgt_5_637;
         Mult_Buf[50].Feature_n = FeatureBuf_638;
         Mult_Buf[50].Weight_n = Wgt_5_638;
         Mult_Buf[51].Feature_n = FeatureBuf_639;
         Mult_Buf[51].Weight_n = Wgt_5_639;
         Mult_Buf[52].Feature_n = FeatureBuf_640;
         Mult_Buf[52].Weight_n = Wgt_5_640;
         Mult_Buf[53].Feature_n = FeatureBuf_641;
         Mult_Buf[53].Weight_n = Wgt_5_641;
         Mult_Buf[54].Feature_n = FeatureBuf_642;
         Mult_Buf[54].Weight_n = Wgt_5_642;
         Mult_Buf[55].Feature_n = FeatureBuf_643;
         Mult_Buf[55].Weight_n = Wgt_5_643;
         Mult_Buf[56].Feature_n = FeatureBuf_644;
         Mult_Buf[56].Weight_n = Wgt_5_644;
         Mult_Buf[57].Feature_n = FeatureBuf_645;
         Mult_Buf[57].Weight_n = Wgt_5_645;
         Mult_Buf[58].Feature_n = FeatureBuf_646;
         Mult_Buf[58].Weight_n = Wgt_5_646;
         Mult_Buf[59].Feature_n = FeatureBuf_647;
         Mult_Buf[59].Weight_n = Wgt_5_647;
         Mult_Buf[60].Feature_n = FeatureBuf_648;
         Mult_Buf[60].Weight_n = Wgt_5_648;
         Mult_Buf[61].Feature_n = FeatureBuf_649;
         Mult_Buf[61].Weight_n = Wgt_5_649;
         Mult_Buf[62].Feature_n = FeatureBuf_650;
         Mult_Buf[62].Weight_n = Wgt_5_650;
         Mult_Buf[63].Feature_n = FeatureBuf_651;
         Mult_Buf[63].Weight_n = Wgt_5_651;
         Mult_Buf[64].Feature_n = FeatureBuf_652;
         Mult_Buf[64].Weight_n = Wgt_5_652;
         Mult_Buf[65].Feature_n = FeatureBuf_653;
         Mult_Buf[65].Weight_n = Wgt_5_653;
         Mult_Buf[66].Feature_n = FeatureBuf_654;
         Mult_Buf[66].Weight_n = Wgt_5_654;
         Mult_Buf[67].Feature_n = FeatureBuf_655;
         Mult_Buf[67].Weight_n = Wgt_5_655;
         Mult_Buf[68].Feature_n = FeatureBuf_656;
         Mult_Buf[68].Weight_n = Wgt_5_656;
         Mult_Buf[69].Feature_n = FeatureBuf_657;
         Mult_Buf[69].Weight_n = Wgt_5_657;
         Mult_Buf[70].Feature_n = FeatureBuf_658;
         Mult_Buf[70].Weight_n = Wgt_5_658;
         Mult_Buf[71].Feature_n = FeatureBuf_659;
         Mult_Buf[71].Weight_n = Wgt_5_659;
         Mult_Buf[72].Feature_n = FeatureBuf_660;
         Mult_Buf[72].Weight_n = Wgt_5_660;
         Mult_Buf[73].Feature_n = FeatureBuf_661;
         Mult_Buf[73].Weight_n = Wgt_5_661;
         Mult_Buf[74].Feature_n = FeatureBuf_662;
         Mult_Buf[74].Weight_n = Wgt_5_662;
         Mult_Buf[75].Feature_n = FeatureBuf_663;
         Mult_Buf[75].Weight_n = Wgt_5_663;
         Mult_Buf[76].Feature_n = FeatureBuf_664;
         Mult_Buf[76].Weight_n = Wgt_5_664;
         Mult_Buf[77].Feature_n = FeatureBuf_665;
         Mult_Buf[77].Weight_n = Wgt_5_665;
         Mult_Buf[78].Feature_n = FeatureBuf_666;
         Mult_Buf[78].Weight_n = Wgt_5_666;
         Mult_Buf[79].Feature_n = FeatureBuf_667;
         Mult_Buf[79].Weight_n = Wgt_5_667;
         Mult_Buf[80].Feature_n = FeatureBuf_668;
         Mult_Buf[80].Weight_n = Wgt_5_668;
         Mult_Buf[81].Feature_n = FeatureBuf_669;
         Mult_Buf[81].Weight_n = Wgt_5_669;
         Mult_Buf[82].Feature_n = FeatureBuf_670;
         Mult_Buf[82].Weight_n = Wgt_5_670;
         Mult_Buf[83].Feature_n = FeatureBuf_671;
         Mult_Buf[83].Weight_n = Wgt_5_671;
         Mult_Buf[84].Feature_n = FeatureBuf_672;
         Mult_Buf[84].Weight_n = Wgt_5_672;
         Mult_Buf[85].Feature_n = FeatureBuf_673;
         Mult_Buf[85].Weight_n = Wgt_5_673;
         Mult_Buf[86].Feature_n = FeatureBuf_674;
         Mult_Buf[86].Weight_n = Wgt_5_674;
         Mult_Buf[87].Feature_n = FeatureBuf_675;
         Mult_Buf[87].Weight_n = Wgt_5_675;
         Mult_Buf[88].Feature_n = FeatureBuf_676;
         Mult_Buf[88].Weight_n = Wgt_5_676;
         Mult_Buf[89].Feature_n = FeatureBuf_677;
         Mult_Buf[89].Weight_n = Wgt_5_677;
         Mult_Buf[90].Feature_n = FeatureBuf_678;
         Mult_Buf[90].Weight_n = Wgt_5_678;
         Mult_Buf[91].Feature_n = FeatureBuf_679;
         Mult_Buf[91].Weight_n = Wgt_5_679;
         Mult_Buf[92].Feature_n = FeatureBuf_680;
         Mult_Buf[92].Weight_n = Wgt_5_680;
         Mult_Buf[93].Feature_n = FeatureBuf_681;
         Mult_Buf[93].Weight_n = Wgt_5_681;
         Mult_Buf[94].Feature_n = FeatureBuf_682;
         Mult_Buf[94].Weight_n = Wgt_5_682;
         Mult_Buf[95].Feature_n = FeatureBuf_683;
         Mult_Buf[95].Weight_n = Wgt_5_683;
         Mult_Buf[96].Feature_n = FeatureBuf_684;
         Mult_Buf[96].Weight_n = Wgt_5_684;
         Mult_Buf[97].Feature_n = FeatureBuf_685;
         Mult_Buf[97].Weight_n = Wgt_5_685;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     //Collect Partial result form Adder
         Res_3_0_n = Part_Res;
     end
    49:begin
     nxt_state = 50;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_686;
         Mult_Buf[0].Weight_n = Wgt_5_686;
         Mult_Buf[1].Feature_n = FeatureBuf_687;
         Mult_Buf[1].Weight_n = Wgt_5_687;
         Mult_Buf[2].Feature_n = FeatureBuf_688;
         Mult_Buf[2].Weight_n = Wgt_5_688;
         Mult_Buf[3].Feature_n = FeatureBuf_689;
         Mult_Buf[3].Weight_n = Wgt_5_689;
         Mult_Buf[4].Feature_n = FeatureBuf_690;
         Mult_Buf[4].Weight_n = Wgt_5_690;
         Mult_Buf[5].Feature_n = FeatureBuf_691;
         Mult_Buf[5].Weight_n = Wgt_5_691;
         Mult_Buf[6].Feature_n = FeatureBuf_692;
         Mult_Buf[6].Weight_n = Wgt_5_692;
         Mult_Buf[7].Feature_n = FeatureBuf_693;
         Mult_Buf[7].Weight_n = Wgt_5_693;
         Mult_Buf[8].Feature_n = FeatureBuf_694;
         Mult_Buf[8].Weight_n = Wgt_5_694;
         Mult_Buf[9].Feature_n = FeatureBuf_695;
         Mult_Buf[9].Weight_n = Wgt_5_695;
         Mult_Buf[10].Feature_n = FeatureBuf_696;
         Mult_Buf[10].Weight_n = Wgt_5_696;
         Mult_Buf[11].Feature_n = FeatureBuf_697;
         Mult_Buf[11].Weight_n = Wgt_5_697;
         Mult_Buf[12].Feature_n = FeatureBuf_698;
         Mult_Buf[12].Weight_n = Wgt_5_698;
         Mult_Buf[13].Feature_n = FeatureBuf_699;
         Mult_Buf[13].Weight_n = Wgt_5_699;
         Mult_Buf[14].Feature_n = FeatureBuf_700;
         Mult_Buf[14].Weight_n = Wgt_5_700;
         Mult_Buf[15].Feature_n = FeatureBuf_701;
         Mult_Buf[15].Weight_n = Wgt_5_701;
         Mult_Buf[16].Feature_n = FeatureBuf_702;
         Mult_Buf[16].Weight_n = Wgt_5_702;
         Mult_Buf[17].Feature_n = FeatureBuf_703;
         Mult_Buf[17].Weight_n = Wgt_5_703;
         Mult_Buf[18].Feature_n = FeatureBuf_704;
         Mult_Buf[18].Weight_n = Wgt_5_704;
         Mult_Buf[19].Feature_n = FeatureBuf_705;
         Mult_Buf[19].Weight_n = Wgt_5_705;
         Mult_Buf[20].Feature_n = FeatureBuf_706;
         Mult_Buf[20].Weight_n = Wgt_5_706;
         Mult_Buf[21].Feature_n = FeatureBuf_707;
         Mult_Buf[21].Weight_n = Wgt_5_707;
         Mult_Buf[22].Feature_n = FeatureBuf_708;
         Mult_Buf[22].Weight_n = Wgt_5_708;
         Mult_Buf[23].Feature_n = FeatureBuf_709;
         Mult_Buf[23].Weight_n = Wgt_5_709;
         Mult_Buf[24].Feature_n = FeatureBuf_710;
         Mult_Buf[24].Weight_n = Wgt_5_710;
         Mult_Buf[25].Feature_n = FeatureBuf_711;
         Mult_Buf[25].Weight_n = Wgt_5_711;
         Mult_Buf[26].Feature_n = FeatureBuf_712;
         Mult_Buf[26].Weight_n = Wgt_5_712;
         Mult_Buf[27].Feature_n = FeatureBuf_713;
         Mult_Buf[27].Weight_n = Wgt_5_713;
         Mult_Buf[28].Feature_n = FeatureBuf_714;
         Mult_Buf[28].Weight_n = Wgt_5_714;
         Mult_Buf[29].Feature_n = FeatureBuf_715;
         Mult_Buf[29].Weight_n = Wgt_5_715;
         Mult_Buf[30].Feature_n = FeatureBuf_716;
         Mult_Buf[30].Weight_n = Wgt_5_716;
         Mult_Buf[31].Feature_n = FeatureBuf_717;
         Mult_Buf[31].Weight_n = Wgt_5_717;
         Mult_Buf[32].Feature_n = FeatureBuf_718;
         Mult_Buf[32].Weight_n = Wgt_5_718;
         Mult_Buf[33].Feature_n = FeatureBuf_719;
         Mult_Buf[33].Weight_n = Wgt_5_719;
         Mult_Buf[34].Feature_n = FeatureBuf_720;
         Mult_Buf[34].Weight_n = Wgt_5_720;
         Mult_Buf[35].Feature_n = FeatureBuf_721;
         Mult_Buf[35].Weight_n = Wgt_5_721;
         Mult_Buf[36].Feature_n = FeatureBuf_722;
         Mult_Buf[36].Weight_n = Wgt_5_722;
         Mult_Buf[37].Feature_n = FeatureBuf_723;
         Mult_Buf[37].Weight_n = Wgt_5_723;
         Mult_Buf[38].Feature_n = FeatureBuf_724;
         Mult_Buf[38].Weight_n = Wgt_5_724;
         Mult_Buf[39].Feature_n = FeatureBuf_725;
         Mult_Buf[39].Weight_n = Wgt_5_725;
         Mult_Buf[40].Feature_n = FeatureBuf_726;
         Mult_Buf[40].Weight_n = Wgt_5_726;
         Mult_Buf[41].Feature_n = FeatureBuf_727;
         Mult_Buf[41].Weight_n = Wgt_5_727;
         Mult_Buf[42].Feature_n = FeatureBuf_728;
         Mult_Buf[42].Weight_n = Wgt_5_728;
         Mult_Buf[43].Feature_n = FeatureBuf_729;
         Mult_Buf[43].Weight_n = Wgt_5_729;
         Mult_Buf[44].Feature_n = FeatureBuf_730;
         Mult_Buf[44].Weight_n = Wgt_5_730;
         Mult_Buf[45].Feature_n = FeatureBuf_731;
         Mult_Buf[45].Weight_n = Wgt_5_731;
         Mult_Buf[46].Feature_n = FeatureBuf_732;
         Mult_Buf[46].Weight_n = Wgt_5_732;
         Mult_Buf[47].Feature_n = FeatureBuf_733;
         Mult_Buf[47].Weight_n = Wgt_5_733;
         Mult_Buf[48].Feature_n = FeatureBuf_734;
         Mult_Buf[48].Weight_n = Wgt_5_734;
         Mult_Buf[49].Feature_n = FeatureBuf_735;
         Mult_Buf[49].Weight_n = Wgt_5_735;
         Mult_Buf[50].Feature_n = FeatureBuf_736;
         Mult_Buf[50].Weight_n = Wgt_5_736;
         Mult_Buf[51].Feature_n = FeatureBuf_737;
         Mult_Buf[51].Weight_n = Wgt_5_737;
         Mult_Buf[52].Feature_n = FeatureBuf_738;
         Mult_Buf[52].Weight_n = Wgt_5_738;
         Mult_Buf[53].Feature_n = FeatureBuf_739;
         Mult_Buf[53].Weight_n = Wgt_5_739;
         Mult_Buf[54].Feature_n = FeatureBuf_740;
         Mult_Buf[54].Weight_n = Wgt_5_740;
         Mult_Buf[55].Feature_n = FeatureBuf_741;
         Mult_Buf[55].Weight_n = Wgt_5_741;
         Mult_Buf[56].Feature_n = FeatureBuf_742;
         Mult_Buf[56].Weight_n = Wgt_5_742;
         Mult_Buf[57].Feature_n = FeatureBuf_743;
         Mult_Buf[57].Weight_n = Wgt_5_743;
         Mult_Buf[58].Feature_n = FeatureBuf_744;
         Mult_Buf[58].Weight_n = Wgt_5_744;
         Mult_Buf[59].Feature_n = FeatureBuf_745;
         Mult_Buf[59].Weight_n = Wgt_5_745;
         Mult_Buf[60].Feature_n = FeatureBuf_746;
         Mult_Buf[60].Weight_n = Wgt_5_746;
         Mult_Buf[61].Feature_n = FeatureBuf_747;
         Mult_Buf[61].Weight_n = Wgt_5_747;
         Mult_Buf[62].Feature_n = FeatureBuf_748;
         Mult_Buf[62].Weight_n = Wgt_5_748;
         Mult_Buf[63].Feature_n = FeatureBuf_749;
         Mult_Buf[63].Weight_n = Wgt_5_749;
         Mult_Buf[64].Feature_n = FeatureBuf_750;
         Mult_Buf[64].Weight_n = Wgt_5_750;
         Mult_Buf[65].Feature_n = FeatureBuf_751;
         Mult_Buf[65].Weight_n = Wgt_5_751;
         Mult_Buf[66].Feature_n = FeatureBuf_752;
         Mult_Buf[66].Weight_n = Wgt_5_752;
         Mult_Buf[67].Feature_n = FeatureBuf_753;
         Mult_Buf[67].Weight_n = Wgt_5_753;
         Mult_Buf[68].Feature_n = FeatureBuf_754;
         Mult_Buf[68].Weight_n = Wgt_5_754;
         Mult_Buf[69].Feature_n = FeatureBuf_755;
         Mult_Buf[69].Weight_n = Wgt_5_755;
         Mult_Buf[70].Feature_n = FeatureBuf_756;
         Mult_Buf[70].Weight_n = Wgt_5_756;
         Mult_Buf[71].Feature_n = FeatureBuf_757;
         Mult_Buf[71].Weight_n = Wgt_5_757;
         Mult_Buf[72].Feature_n = FeatureBuf_758;
         Mult_Buf[72].Weight_n = Wgt_5_758;
         Mult_Buf[73].Feature_n = FeatureBuf_759;
         Mult_Buf[73].Weight_n = Wgt_5_759;
         Mult_Buf[74].Feature_n = FeatureBuf_760;
         Mult_Buf[74].Weight_n = Wgt_5_760;
         Mult_Buf[75].Feature_n = FeatureBuf_761;
         Mult_Buf[75].Weight_n = Wgt_5_761;
         Mult_Buf[76].Feature_n = FeatureBuf_762;
         Mult_Buf[76].Weight_n = Wgt_5_762;
         Mult_Buf[77].Feature_n = FeatureBuf_763;
         Mult_Buf[77].Weight_n = Wgt_5_763;
         Mult_Buf[78].Feature_n = FeatureBuf_764;
         Mult_Buf[78].Weight_n = Wgt_5_764;
         Mult_Buf[79].Feature_n = FeatureBuf_765;
         Mult_Buf[79].Weight_n = Wgt_5_765;
         Mult_Buf[80].Feature_n = FeatureBuf_766;
         Mult_Buf[80].Weight_n = Wgt_5_766;
         Mult_Buf[81].Feature_n = FeatureBuf_767;
         Mult_Buf[81].Weight_n = Wgt_5_767;
         Mult_Buf[82].Feature_n = FeatureBuf_768;
         Mult_Buf[82].Weight_n = Wgt_5_768;
         Mult_Buf[83].Feature_n = FeatureBuf_769;
         Mult_Buf[83].Weight_n = Wgt_5_769;
         Mult_Buf[84].Feature_n = FeatureBuf_770;
         Mult_Buf[84].Weight_n = Wgt_5_770;
         Mult_Buf[85].Feature_n = FeatureBuf_771;
         Mult_Buf[85].Weight_n = Wgt_5_771;
         Mult_Buf[86].Feature_n = FeatureBuf_772;
         Mult_Buf[86].Weight_n = Wgt_5_772;
         Mult_Buf[87].Feature_n = FeatureBuf_773;
         Mult_Buf[87].Weight_n = Wgt_5_773;
         Mult_Buf[88].Feature_n = FeatureBuf_774;
         Mult_Buf[88].Weight_n = Wgt_5_774;
         Mult_Buf[89].Feature_n = FeatureBuf_775;
         Mult_Buf[89].Weight_n = Wgt_5_775;
         Mult_Buf[90].Feature_n = FeatureBuf_776;
         Mult_Buf[90].Weight_n = Wgt_5_776;
         Mult_Buf[91].Feature_n = FeatureBuf_777;
         Mult_Buf[91].Weight_n = Wgt_5_777;
         Mult_Buf[92].Feature_n = FeatureBuf_778;
         Mult_Buf[92].Weight_n = Wgt_5_778;
         Mult_Buf[93].Feature_n = FeatureBuf_779;
         Mult_Buf[93].Weight_n = Wgt_5_779;
         Mult_Buf[94].Feature_n = FeatureBuf_780;
         Mult_Buf[94].Weight_n = Wgt_5_780;
         Mult_Buf[95].Feature_n = FeatureBuf_781;
         Mult_Buf[95].Weight_n = Wgt_5_781;
         Mult_Buf[96].Feature_n = FeatureBuf_782;
         Mult_Buf[96].Weight_n = Wgt_5_782;
         Mult_Buf[97].Feature_n = FeatureBuf_783;
         Mult_Buf[97].Weight_n = Wgt_5_783;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     //Collect Partial result form Adder
         Res_3_1_n = Part_Res;
     end
    50:begin
     nxt_state = 51;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_0;
         Mult_Buf[0].Weight_n = Wgt_6_0;
         Mult_Buf[1].Feature_n = FeatureBuf_1;
         Mult_Buf[1].Weight_n = Wgt_6_1;
         Mult_Buf[2].Feature_n = FeatureBuf_2;
         Mult_Buf[2].Weight_n = Wgt_6_2;
         Mult_Buf[3].Feature_n = FeatureBuf_3;
         Mult_Buf[3].Weight_n = Wgt_6_3;
         Mult_Buf[4].Feature_n = FeatureBuf_4;
         Mult_Buf[4].Weight_n = Wgt_6_4;
         Mult_Buf[5].Feature_n = FeatureBuf_5;
         Mult_Buf[5].Weight_n = Wgt_6_5;
         Mult_Buf[6].Feature_n = FeatureBuf_6;
         Mult_Buf[6].Weight_n = Wgt_6_6;
         Mult_Buf[7].Feature_n = FeatureBuf_7;
         Mult_Buf[7].Weight_n = Wgt_6_7;
         Mult_Buf[8].Feature_n = FeatureBuf_8;
         Mult_Buf[8].Weight_n = Wgt_6_8;
         Mult_Buf[9].Feature_n = FeatureBuf_9;
         Mult_Buf[9].Weight_n = Wgt_6_9;
         Mult_Buf[10].Feature_n = FeatureBuf_10;
         Mult_Buf[10].Weight_n = Wgt_6_10;
         Mult_Buf[11].Feature_n = FeatureBuf_11;
         Mult_Buf[11].Weight_n = Wgt_6_11;
         Mult_Buf[12].Feature_n = FeatureBuf_12;
         Mult_Buf[12].Weight_n = Wgt_6_12;
         Mult_Buf[13].Feature_n = FeatureBuf_13;
         Mult_Buf[13].Weight_n = Wgt_6_13;
         Mult_Buf[14].Feature_n = FeatureBuf_14;
         Mult_Buf[14].Weight_n = Wgt_6_14;
         Mult_Buf[15].Feature_n = FeatureBuf_15;
         Mult_Buf[15].Weight_n = Wgt_6_15;
         Mult_Buf[16].Feature_n = FeatureBuf_16;
         Mult_Buf[16].Weight_n = Wgt_6_16;
         Mult_Buf[17].Feature_n = FeatureBuf_17;
         Mult_Buf[17].Weight_n = Wgt_6_17;
         Mult_Buf[18].Feature_n = FeatureBuf_18;
         Mult_Buf[18].Weight_n = Wgt_6_18;
         Mult_Buf[19].Feature_n = FeatureBuf_19;
         Mult_Buf[19].Weight_n = Wgt_6_19;
         Mult_Buf[20].Feature_n = FeatureBuf_20;
         Mult_Buf[20].Weight_n = Wgt_6_20;
         Mult_Buf[21].Feature_n = FeatureBuf_21;
         Mult_Buf[21].Weight_n = Wgt_6_21;
         Mult_Buf[22].Feature_n = FeatureBuf_22;
         Mult_Buf[22].Weight_n = Wgt_6_22;
         Mult_Buf[23].Feature_n = FeatureBuf_23;
         Mult_Buf[23].Weight_n = Wgt_6_23;
         Mult_Buf[24].Feature_n = FeatureBuf_24;
         Mult_Buf[24].Weight_n = Wgt_6_24;
         Mult_Buf[25].Feature_n = FeatureBuf_25;
         Mult_Buf[25].Weight_n = Wgt_6_25;
         Mult_Buf[26].Feature_n = FeatureBuf_26;
         Mult_Buf[26].Weight_n = Wgt_6_26;
         Mult_Buf[27].Feature_n = FeatureBuf_27;
         Mult_Buf[27].Weight_n = Wgt_6_27;
         Mult_Buf[28].Feature_n = FeatureBuf_28;
         Mult_Buf[28].Weight_n = Wgt_6_28;
         Mult_Buf[29].Feature_n = FeatureBuf_29;
         Mult_Buf[29].Weight_n = Wgt_6_29;
         Mult_Buf[30].Feature_n = FeatureBuf_30;
         Mult_Buf[30].Weight_n = Wgt_6_30;
         Mult_Buf[31].Feature_n = FeatureBuf_31;
         Mult_Buf[31].Weight_n = Wgt_6_31;
         Mult_Buf[32].Feature_n = FeatureBuf_32;
         Mult_Buf[32].Weight_n = Wgt_6_32;
         Mult_Buf[33].Feature_n = FeatureBuf_33;
         Mult_Buf[33].Weight_n = Wgt_6_33;
         Mult_Buf[34].Feature_n = FeatureBuf_34;
         Mult_Buf[34].Weight_n = Wgt_6_34;
         Mult_Buf[35].Feature_n = FeatureBuf_35;
         Mult_Buf[35].Weight_n = Wgt_6_35;
         Mult_Buf[36].Feature_n = FeatureBuf_36;
         Mult_Buf[36].Weight_n = Wgt_6_36;
         Mult_Buf[37].Feature_n = FeatureBuf_37;
         Mult_Buf[37].Weight_n = Wgt_6_37;
         Mult_Buf[38].Feature_n = FeatureBuf_38;
         Mult_Buf[38].Weight_n = Wgt_6_38;
         Mult_Buf[39].Feature_n = FeatureBuf_39;
         Mult_Buf[39].Weight_n = Wgt_6_39;
         Mult_Buf[40].Feature_n = FeatureBuf_40;
         Mult_Buf[40].Weight_n = Wgt_6_40;
         Mult_Buf[41].Feature_n = FeatureBuf_41;
         Mult_Buf[41].Weight_n = Wgt_6_41;
         Mult_Buf[42].Feature_n = FeatureBuf_42;
         Mult_Buf[42].Weight_n = Wgt_6_42;
         Mult_Buf[43].Feature_n = FeatureBuf_43;
         Mult_Buf[43].Weight_n = Wgt_6_43;
         Mult_Buf[44].Feature_n = FeatureBuf_44;
         Mult_Buf[44].Weight_n = Wgt_6_44;
         Mult_Buf[45].Feature_n = FeatureBuf_45;
         Mult_Buf[45].Weight_n = Wgt_6_45;
         Mult_Buf[46].Feature_n = FeatureBuf_46;
         Mult_Buf[46].Weight_n = Wgt_6_46;
         Mult_Buf[47].Feature_n = FeatureBuf_47;
         Mult_Buf[47].Weight_n = Wgt_6_47;
         Mult_Buf[48].Feature_n = FeatureBuf_48;
         Mult_Buf[48].Weight_n = Wgt_6_48;
         Mult_Buf[49].Feature_n = FeatureBuf_49;
         Mult_Buf[49].Weight_n = Wgt_6_49;
         Mult_Buf[50].Feature_n = FeatureBuf_50;
         Mult_Buf[50].Weight_n = Wgt_6_50;
         Mult_Buf[51].Feature_n = FeatureBuf_51;
         Mult_Buf[51].Weight_n = Wgt_6_51;
         Mult_Buf[52].Feature_n = FeatureBuf_52;
         Mult_Buf[52].Weight_n = Wgt_6_52;
         Mult_Buf[53].Feature_n = FeatureBuf_53;
         Mult_Buf[53].Weight_n = Wgt_6_53;
         Mult_Buf[54].Feature_n = FeatureBuf_54;
         Mult_Buf[54].Weight_n = Wgt_6_54;
         Mult_Buf[55].Feature_n = FeatureBuf_55;
         Mult_Buf[55].Weight_n = Wgt_6_55;
         Mult_Buf[56].Feature_n = FeatureBuf_56;
         Mult_Buf[56].Weight_n = Wgt_6_56;
         Mult_Buf[57].Feature_n = FeatureBuf_57;
         Mult_Buf[57].Weight_n = Wgt_6_57;
         Mult_Buf[58].Feature_n = FeatureBuf_58;
         Mult_Buf[58].Weight_n = Wgt_6_58;
         Mult_Buf[59].Feature_n = FeatureBuf_59;
         Mult_Buf[59].Weight_n = Wgt_6_59;
         Mult_Buf[60].Feature_n = FeatureBuf_60;
         Mult_Buf[60].Weight_n = Wgt_6_60;
         Mult_Buf[61].Feature_n = FeatureBuf_61;
         Mult_Buf[61].Weight_n = Wgt_6_61;
         Mult_Buf[62].Feature_n = FeatureBuf_62;
         Mult_Buf[62].Weight_n = Wgt_6_62;
         Mult_Buf[63].Feature_n = FeatureBuf_63;
         Mult_Buf[63].Weight_n = Wgt_6_63;
         Mult_Buf[64].Feature_n = FeatureBuf_64;
         Mult_Buf[64].Weight_n = Wgt_6_64;
         Mult_Buf[65].Feature_n = FeatureBuf_65;
         Mult_Buf[65].Weight_n = Wgt_6_65;
         Mult_Buf[66].Feature_n = FeatureBuf_66;
         Mult_Buf[66].Weight_n = Wgt_6_66;
         Mult_Buf[67].Feature_n = FeatureBuf_67;
         Mult_Buf[67].Weight_n = Wgt_6_67;
         Mult_Buf[68].Feature_n = FeatureBuf_68;
         Mult_Buf[68].Weight_n = Wgt_6_68;
         Mult_Buf[69].Feature_n = FeatureBuf_69;
         Mult_Buf[69].Weight_n = Wgt_6_69;
         Mult_Buf[70].Feature_n = FeatureBuf_70;
         Mult_Buf[70].Weight_n = Wgt_6_70;
         Mult_Buf[71].Feature_n = FeatureBuf_71;
         Mult_Buf[71].Weight_n = Wgt_6_71;
         Mult_Buf[72].Feature_n = FeatureBuf_72;
         Mult_Buf[72].Weight_n = Wgt_6_72;
         Mult_Buf[73].Feature_n = FeatureBuf_73;
         Mult_Buf[73].Weight_n = Wgt_6_73;
         Mult_Buf[74].Feature_n = FeatureBuf_74;
         Mult_Buf[74].Weight_n = Wgt_6_74;
         Mult_Buf[75].Feature_n = FeatureBuf_75;
         Mult_Buf[75].Weight_n = Wgt_6_75;
         Mult_Buf[76].Feature_n = FeatureBuf_76;
         Mult_Buf[76].Weight_n = Wgt_6_76;
         Mult_Buf[77].Feature_n = FeatureBuf_77;
         Mult_Buf[77].Weight_n = Wgt_6_77;
         Mult_Buf[78].Feature_n = FeatureBuf_78;
         Mult_Buf[78].Weight_n = Wgt_6_78;
         Mult_Buf[79].Feature_n = FeatureBuf_79;
         Mult_Buf[79].Weight_n = Wgt_6_79;
         Mult_Buf[80].Feature_n = FeatureBuf_80;
         Mult_Buf[80].Weight_n = Wgt_6_80;
         Mult_Buf[81].Feature_n = FeatureBuf_81;
         Mult_Buf[81].Weight_n = Wgt_6_81;
         Mult_Buf[82].Feature_n = FeatureBuf_82;
         Mult_Buf[82].Weight_n = Wgt_6_82;
         Mult_Buf[83].Feature_n = FeatureBuf_83;
         Mult_Buf[83].Weight_n = Wgt_6_83;
         Mult_Buf[84].Feature_n = FeatureBuf_84;
         Mult_Buf[84].Weight_n = Wgt_6_84;
         Mult_Buf[85].Feature_n = FeatureBuf_85;
         Mult_Buf[85].Weight_n = Wgt_6_85;
         Mult_Buf[86].Feature_n = FeatureBuf_86;
         Mult_Buf[86].Weight_n = Wgt_6_86;
         Mult_Buf[87].Feature_n = FeatureBuf_87;
         Mult_Buf[87].Weight_n = Wgt_6_87;
         Mult_Buf[88].Feature_n = FeatureBuf_88;
         Mult_Buf[88].Weight_n = Wgt_6_88;
         Mult_Buf[89].Feature_n = FeatureBuf_89;
         Mult_Buf[89].Weight_n = Wgt_6_89;
         Mult_Buf[90].Feature_n = FeatureBuf_90;
         Mult_Buf[90].Weight_n = Wgt_6_90;
         Mult_Buf[91].Feature_n = FeatureBuf_91;
         Mult_Buf[91].Weight_n = Wgt_6_91;
         Mult_Buf[92].Feature_n = FeatureBuf_92;
         Mult_Buf[92].Weight_n = Wgt_6_92;
         Mult_Buf[93].Feature_n = FeatureBuf_93;
         Mult_Buf[93].Weight_n = Wgt_6_93;
         Mult_Buf[94].Feature_n = FeatureBuf_94;
         Mult_Buf[94].Weight_n = Wgt_6_94;
         Mult_Buf[95].Feature_n = FeatureBuf_95;
         Mult_Buf[95].Weight_n = Wgt_6_95;
         Mult_Buf[96].Feature_n = FeatureBuf_96;
         Mult_Buf[96].Weight_n = Wgt_6_96;
         Mult_Buf[97].Feature_n = FeatureBuf_97;
         Mult_Buf[97].Weight_n = Wgt_6_97;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     //Collect Partial result form Adder
         Res_3_2_n = Part_Res;
     end
    51:begin
     nxt_state = 52;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_98;
         Mult_Buf[0].Weight_n = Wgt_6_98;
         Mult_Buf[1].Feature_n = FeatureBuf_99;
         Mult_Buf[1].Weight_n = Wgt_6_99;
         Mult_Buf[2].Feature_n = FeatureBuf_100;
         Mult_Buf[2].Weight_n = Wgt_6_100;
         Mult_Buf[3].Feature_n = FeatureBuf_101;
         Mult_Buf[3].Weight_n = Wgt_6_101;
         Mult_Buf[4].Feature_n = FeatureBuf_102;
         Mult_Buf[4].Weight_n = Wgt_6_102;
         Mult_Buf[5].Feature_n = FeatureBuf_103;
         Mult_Buf[5].Weight_n = Wgt_6_103;
         Mult_Buf[6].Feature_n = FeatureBuf_104;
         Mult_Buf[6].Weight_n = Wgt_6_104;
         Mult_Buf[7].Feature_n = FeatureBuf_105;
         Mult_Buf[7].Weight_n = Wgt_6_105;
         Mult_Buf[8].Feature_n = FeatureBuf_106;
         Mult_Buf[8].Weight_n = Wgt_6_106;
         Mult_Buf[9].Feature_n = FeatureBuf_107;
         Mult_Buf[9].Weight_n = Wgt_6_107;
         Mult_Buf[10].Feature_n = FeatureBuf_108;
         Mult_Buf[10].Weight_n = Wgt_6_108;
         Mult_Buf[11].Feature_n = FeatureBuf_109;
         Mult_Buf[11].Weight_n = Wgt_6_109;
         Mult_Buf[12].Feature_n = FeatureBuf_110;
         Mult_Buf[12].Weight_n = Wgt_6_110;
         Mult_Buf[13].Feature_n = FeatureBuf_111;
         Mult_Buf[13].Weight_n = Wgt_6_111;
         Mult_Buf[14].Feature_n = FeatureBuf_112;
         Mult_Buf[14].Weight_n = Wgt_6_112;
         Mult_Buf[15].Feature_n = FeatureBuf_113;
         Mult_Buf[15].Weight_n = Wgt_6_113;
         Mult_Buf[16].Feature_n = FeatureBuf_114;
         Mult_Buf[16].Weight_n = Wgt_6_114;
         Mult_Buf[17].Feature_n = FeatureBuf_115;
         Mult_Buf[17].Weight_n = Wgt_6_115;
         Mult_Buf[18].Feature_n = FeatureBuf_116;
         Mult_Buf[18].Weight_n = Wgt_6_116;
         Mult_Buf[19].Feature_n = FeatureBuf_117;
         Mult_Buf[19].Weight_n = Wgt_6_117;
         Mult_Buf[20].Feature_n = FeatureBuf_118;
         Mult_Buf[20].Weight_n = Wgt_6_118;
         Mult_Buf[21].Feature_n = FeatureBuf_119;
         Mult_Buf[21].Weight_n = Wgt_6_119;
         Mult_Buf[22].Feature_n = FeatureBuf_120;
         Mult_Buf[22].Weight_n = Wgt_6_120;
         Mult_Buf[23].Feature_n = FeatureBuf_121;
         Mult_Buf[23].Weight_n = Wgt_6_121;
         Mult_Buf[24].Feature_n = FeatureBuf_122;
         Mult_Buf[24].Weight_n = Wgt_6_122;
         Mult_Buf[25].Feature_n = FeatureBuf_123;
         Mult_Buf[25].Weight_n = Wgt_6_123;
         Mult_Buf[26].Feature_n = FeatureBuf_124;
         Mult_Buf[26].Weight_n = Wgt_6_124;
         Mult_Buf[27].Feature_n = FeatureBuf_125;
         Mult_Buf[27].Weight_n = Wgt_6_125;
         Mult_Buf[28].Feature_n = FeatureBuf_126;
         Mult_Buf[28].Weight_n = Wgt_6_126;
         Mult_Buf[29].Feature_n = FeatureBuf_127;
         Mult_Buf[29].Weight_n = Wgt_6_127;
         Mult_Buf[30].Feature_n = FeatureBuf_128;
         Mult_Buf[30].Weight_n = Wgt_6_128;
         Mult_Buf[31].Feature_n = FeatureBuf_129;
         Mult_Buf[31].Weight_n = Wgt_6_129;
         Mult_Buf[32].Feature_n = FeatureBuf_130;
         Mult_Buf[32].Weight_n = Wgt_6_130;
         Mult_Buf[33].Feature_n = FeatureBuf_131;
         Mult_Buf[33].Weight_n = Wgt_6_131;
         Mult_Buf[34].Feature_n = FeatureBuf_132;
         Mult_Buf[34].Weight_n = Wgt_6_132;
         Mult_Buf[35].Feature_n = FeatureBuf_133;
         Mult_Buf[35].Weight_n = Wgt_6_133;
         Mult_Buf[36].Feature_n = FeatureBuf_134;
         Mult_Buf[36].Weight_n = Wgt_6_134;
         Mult_Buf[37].Feature_n = FeatureBuf_135;
         Mult_Buf[37].Weight_n = Wgt_6_135;
         Mult_Buf[38].Feature_n = FeatureBuf_136;
         Mult_Buf[38].Weight_n = Wgt_6_136;
         Mult_Buf[39].Feature_n = FeatureBuf_137;
         Mult_Buf[39].Weight_n = Wgt_6_137;
         Mult_Buf[40].Feature_n = FeatureBuf_138;
         Mult_Buf[40].Weight_n = Wgt_6_138;
         Mult_Buf[41].Feature_n = FeatureBuf_139;
         Mult_Buf[41].Weight_n = Wgt_6_139;
         Mult_Buf[42].Feature_n = FeatureBuf_140;
         Mult_Buf[42].Weight_n = Wgt_6_140;
         Mult_Buf[43].Feature_n = FeatureBuf_141;
         Mult_Buf[43].Weight_n = Wgt_6_141;
         Mult_Buf[44].Feature_n = FeatureBuf_142;
         Mult_Buf[44].Weight_n = Wgt_6_142;
         Mult_Buf[45].Feature_n = FeatureBuf_143;
         Mult_Buf[45].Weight_n = Wgt_6_143;
         Mult_Buf[46].Feature_n = FeatureBuf_144;
         Mult_Buf[46].Weight_n = Wgt_6_144;
         Mult_Buf[47].Feature_n = FeatureBuf_145;
         Mult_Buf[47].Weight_n = Wgt_6_145;
         Mult_Buf[48].Feature_n = FeatureBuf_146;
         Mult_Buf[48].Weight_n = Wgt_6_146;
         Mult_Buf[49].Feature_n = FeatureBuf_147;
         Mult_Buf[49].Weight_n = Wgt_6_147;
         Mult_Buf[50].Feature_n = FeatureBuf_148;
         Mult_Buf[50].Weight_n = Wgt_6_148;
         Mult_Buf[51].Feature_n = FeatureBuf_149;
         Mult_Buf[51].Weight_n = Wgt_6_149;
         Mult_Buf[52].Feature_n = FeatureBuf_150;
         Mult_Buf[52].Weight_n = Wgt_6_150;
         Mult_Buf[53].Feature_n = FeatureBuf_151;
         Mult_Buf[53].Weight_n = Wgt_6_151;
         Mult_Buf[54].Feature_n = FeatureBuf_152;
         Mult_Buf[54].Weight_n = Wgt_6_152;
         Mult_Buf[55].Feature_n = FeatureBuf_153;
         Mult_Buf[55].Weight_n = Wgt_6_153;
         Mult_Buf[56].Feature_n = FeatureBuf_154;
         Mult_Buf[56].Weight_n = Wgt_6_154;
         Mult_Buf[57].Feature_n = FeatureBuf_155;
         Mult_Buf[57].Weight_n = Wgt_6_155;
         Mult_Buf[58].Feature_n = FeatureBuf_156;
         Mult_Buf[58].Weight_n = Wgt_6_156;
         Mult_Buf[59].Feature_n = FeatureBuf_157;
         Mult_Buf[59].Weight_n = Wgt_6_157;
         Mult_Buf[60].Feature_n = FeatureBuf_158;
         Mult_Buf[60].Weight_n = Wgt_6_158;
         Mult_Buf[61].Feature_n = FeatureBuf_159;
         Mult_Buf[61].Weight_n = Wgt_6_159;
         Mult_Buf[62].Feature_n = FeatureBuf_160;
         Mult_Buf[62].Weight_n = Wgt_6_160;
         Mult_Buf[63].Feature_n = FeatureBuf_161;
         Mult_Buf[63].Weight_n = Wgt_6_161;
         Mult_Buf[64].Feature_n = FeatureBuf_162;
         Mult_Buf[64].Weight_n = Wgt_6_162;
         Mult_Buf[65].Feature_n = FeatureBuf_163;
         Mult_Buf[65].Weight_n = Wgt_6_163;
         Mult_Buf[66].Feature_n = FeatureBuf_164;
         Mult_Buf[66].Weight_n = Wgt_6_164;
         Mult_Buf[67].Feature_n = FeatureBuf_165;
         Mult_Buf[67].Weight_n = Wgt_6_165;
         Mult_Buf[68].Feature_n = FeatureBuf_166;
         Mult_Buf[68].Weight_n = Wgt_6_166;
         Mult_Buf[69].Feature_n = FeatureBuf_167;
         Mult_Buf[69].Weight_n = Wgt_6_167;
         Mult_Buf[70].Feature_n = FeatureBuf_168;
         Mult_Buf[70].Weight_n = Wgt_6_168;
         Mult_Buf[71].Feature_n = FeatureBuf_169;
         Mult_Buf[71].Weight_n = Wgt_6_169;
         Mult_Buf[72].Feature_n = FeatureBuf_170;
         Mult_Buf[72].Weight_n = Wgt_6_170;
         Mult_Buf[73].Feature_n = FeatureBuf_171;
         Mult_Buf[73].Weight_n = Wgt_6_171;
         Mult_Buf[74].Feature_n = FeatureBuf_172;
         Mult_Buf[74].Weight_n = Wgt_6_172;
         Mult_Buf[75].Feature_n = FeatureBuf_173;
         Mult_Buf[75].Weight_n = Wgt_6_173;
         Mult_Buf[76].Feature_n = FeatureBuf_174;
         Mult_Buf[76].Weight_n = Wgt_6_174;
         Mult_Buf[77].Feature_n = FeatureBuf_175;
         Mult_Buf[77].Weight_n = Wgt_6_175;
         Mult_Buf[78].Feature_n = FeatureBuf_176;
         Mult_Buf[78].Weight_n = Wgt_6_176;
         Mult_Buf[79].Feature_n = FeatureBuf_177;
         Mult_Buf[79].Weight_n = Wgt_6_177;
         Mult_Buf[80].Feature_n = FeatureBuf_178;
         Mult_Buf[80].Weight_n = Wgt_6_178;
         Mult_Buf[81].Feature_n = FeatureBuf_179;
         Mult_Buf[81].Weight_n = Wgt_6_179;
         Mult_Buf[82].Feature_n = FeatureBuf_180;
         Mult_Buf[82].Weight_n = Wgt_6_180;
         Mult_Buf[83].Feature_n = FeatureBuf_181;
         Mult_Buf[83].Weight_n = Wgt_6_181;
         Mult_Buf[84].Feature_n = FeatureBuf_182;
         Mult_Buf[84].Weight_n = Wgt_6_182;
         Mult_Buf[85].Feature_n = FeatureBuf_183;
         Mult_Buf[85].Weight_n = Wgt_6_183;
         Mult_Buf[86].Feature_n = FeatureBuf_184;
         Mult_Buf[86].Weight_n = Wgt_6_184;
         Mult_Buf[87].Feature_n = FeatureBuf_185;
         Mult_Buf[87].Weight_n = Wgt_6_185;
         Mult_Buf[88].Feature_n = FeatureBuf_186;
         Mult_Buf[88].Weight_n = Wgt_6_186;
         Mult_Buf[89].Feature_n = FeatureBuf_187;
         Mult_Buf[89].Weight_n = Wgt_6_187;
         Mult_Buf[90].Feature_n = FeatureBuf_188;
         Mult_Buf[90].Weight_n = Wgt_6_188;
         Mult_Buf[91].Feature_n = FeatureBuf_189;
         Mult_Buf[91].Weight_n = Wgt_6_189;
         Mult_Buf[92].Feature_n = FeatureBuf_190;
         Mult_Buf[92].Weight_n = Wgt_6_190;
         Mult_Buf[93].Feature_n = FeatureBuf_191;
         Mult_Buf[93].Weight_n = Wgt_6_191;
         Mult_Buf[94].Feature_n = FeatureBuf_192;
         Mult_Buf[94].Weight_n = Wgt_6_192;
         Mult_Buf[95].Feature_n = FeatureBuf_193;
         Mult_Buf[95].Weight_n = Wgt_6_193;
         Mult_Buf[96].Feature_n = FeatureBuf_194;
         Mult_Buf[96].Weight_n = Wgt_6_194;
         Mult_Buf[97].Feature_n = FeatureBuf_195;
         Mult_Buf[97].Weight_n = Wgt_6_195;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     //Collect Partial result form Adder
         Res_3_3_n = Part_Res;
     end
    52:begin
     nxt_state = 53;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_196;
         Mult_Buf[0].Weight_n = Wgt_6_196;
         Mult_Buf[1].Feature_n = FeatureBuf_197;
         Mult_Buf[1].Weight_n = Wgt_6_197;
         Mult_Buf[2].Feature_n = FeatureBuf_198;
         Mult_Buf[2].Weight_n = Wgt_6_198;
         Mult_Buf[3].Feature_n = FeatureBuf_199;
         Mult_Buf[3].Weight_n = Wgt_6_199;
         Mult_Buf[4].Feature_n = FeatureBuf_200;
         Mult_Buf[4].Weight_n = Wgt_6_200;
         Mult_Buf[5].Feature_n = FeatureBuf_201;
         Mult_Buf[5].Weight_n = Wgt_6_201;
         Mult_Buf[6].Feature_n = FeatureBuf_202;
         Mult_Buf[6].Weight_n = Wgt_6_202;
         Mult_Buf[7].Feature_n = FeatureBuf_203;
         Mult_Buf[7].Weight_n = Wgt_6_203;
         Mult_Buf[8].Feature_n = FeatureBuf_204;
         Mult_Buf[8].Weight_n = Wgt_6_204;
         Mult_Buf[9].Feature_n = FeatureBuf_205;
         Mult_Buf[9].Weight_n = Wgt_6_205;
         Mult_Buf[10].Feature_n = FeatureBuf_206;
         Mult_Buf[10].Weight_n = Wgt_6_206;
         Mult_Buf[11].Feature_n = FeatureBuf_207;
         Mult_Buf[11].Weight_n = Wgt_6_207;
         Mult_Buf[12].Feature_n = FeatureBuf_208;
         Mult_Buf[12].Weight_n = Wgt_6_208;
         Mult_Buf[13].Feature_n = FeatureBuf_209;
         Mult_Buf[13].Weight_n = Wgt_6_209;
         Mult_Buf[14].Feature_n = FeatureBuf_210;
         Mult_Buf[14].Weight_n = Wgt_6_210;
         Mult_Buf[15].Feature_n = FeatureBuf_211;
         Mult_Buf[15].Weight_n = Wgt_6_211;
         Mult_Buf[16].Feature_n = FeatureBuf_212;
         Mult_Buf[16].Weight_n = Wgt_6_212;
         Mult_Buf[17].Feature_n = FeatureBuf_213;
         Mult_Buf[17].Weight_n = Wgt_6_213;
         Mult_Buf[18].Feature_n = FeatureBuf_214;
         Mult_Buf[18].Weight_n = Wgt_6_214;
         Mult_Buf[19].Feature_n = FeatureBuf_215;
         Mult_Buf[19].Weight_n = Wgt_6_215;
         Mult_Buf[20].Feature_n = FeatureBuf_216;
         Mult_Buf[20].Weight_n = Wgt_6_216;
         Mult_Buf[21].Feature_n = FeatureBuf_217;
         Mult_Buf[21].Weight_n = Wgt_6_217;
         Mult_Buf[22].Feature_n = FeatureBuf_218;
         Mult_Buf[22].Weight_n = Wgt_6_218;
         Mult_Buf[23].Feature_n = FeatureBuf_219;
         Mult_Buf[23].Weight_n = Wgt_6_219;
         Mult_Buf[24].Feature_n = FeatureBuf_220;
         Mult_Buf[24].Weight_n = Wgt_6_220;
         Mult_Buf[25].Feature_n = FeatureBuf_221;
         Mult_Buf[25].Weight_n = Wgt_6_221;
         Mult_Buf[26].Feature_n = FeatureBuf_222;
         Mult_Buf[26].Weight_n = Wgt_6_222;
         Mult_Buf[27].Feature_n = FeatureBuf_223;
         Mult_Buf[27].Weight_n = Wgt_6_223;
         Mult_Buf[28].Feature_n = FeatureBuf_224;
         Mult_Buf[28].Weight_n = Wgt_6_224;
         Mult_Buf[29].Feature_n = FeatureBuf_225;
         Mult_Buf[29].Weight_n = Wgt_6_225;
         Mult_Buf[30].Feature_n = FeatureBuf_226;
         Mult_Buf[30].Weight_n = Wgt_6_226;
         Mult_Buf[31].Feature_n = FeatureBuf_227;
         Mult_Buf[31].Weight_n = Wgt_6_227;
         Mult_Buf[32].Feature_n = FeatureBuf_228;
         Mult_Buf[32].Weight_n = Wgt_6_228;
         Mult_Buf[33].Feature_n = FeatureBuf_229;
         Mult_Buf[33].Weight_n = Wgt_6_229;
         Mult_Buf[34].Feature_n = FeatureBuf_230;
         Mult_Buf[34].Weight_n = Wgt_6_230;
         Mult_Buf[35].Feature_n = FeatureBuf_231;
         Mult_Buf[35].Weight_n = Wgt_6_231;
         Mult_Buf[36].Feature_n = FeatureBuf_232;
         Mult_Buf[36].Weight_n = Wgt_6_232;
         Mult_Buf[37].Feature_n = FeatureBuf_233;
         Mult_Buf[37].Weight_n = Wgt_6_233;
         Mult_Buf[38].Feature_n = FeatureBuf_234;
         Mult_Buf[38].Weight_n = Wgt_6_234;
         Mult_Buf[39].Feature_n = FeatureBuf_235;
         Mult_Buf[39].Weight_n = Wgt_6_235;
         Mult_Buf[40].Feature_n = FeatureBuf_236;
         Mult_Buf[40].Weight_n = Wgt_6_236;
         Mult_Buf[41].Feature_n = FeatureBuf_237;
         Mult_Buf[41].Weight_n = Wgt_6_237;
         Mult_Buf[42].Feature_n = FeatureBuf_238;
         Mult_Buf[42].Weight_n = Wgt_6_238;
         Mult_Buf[43].Feature_n = FeatureBuf_239;
         Mult_Buf[43].Weight_n = Wgt_6_239;
         Mult_Buf[44].Feature_n = FeatureBuf_240;
         Mult_Buf[44].Weight_n = Wgt_6_240;
         Mult_Buf[45].Feature_n = FeatureBuf_241;
         Mult_Buf[45].Weight_n = Wgt_6_241;
         Mult_Buf[46].Feature_n = FeatureBuf_242;
         Mult_Buf[46].Weight_n = Wgt_6_242;
         Mult_Buf[47].Feature_n = FeatureBuf_243;
         Mult_Buf[47].Weight_n = Wgt_6_243;
         Mult_Buf[48].Feature_n = FeatureBuf_244;
         Mult_Buf[48].Weight_n = Wgt_6_244;
         Mult_Buf[49].Feature_n = FeatureBuf_245;
         Mult_Buf[49].Weight_n = Wgt_6_245;
         Mult_Buf[50].Feature_n = FeatureBuf_246;
         Mult_Buf[50].Weight_n = Wgt_6_246;
         Mult_Buf[51].Feature_n = FeatureBuf_247;
         Mult_Buf[51].Weight_n = Wgt_6_247;
         Mult_Buf[52].Feature_n = FeatureBuf_248;
         Mult_Buf[52].Weight_n = Wgt_6_248;
         Mult_Buf[53].Feature_n = FeatureBuf_249;
         Mult_Buf[53].Weight_n = Wgt_6_249;
         Mult_Buf[54].Feature_n = FeatureBuf_250;
         Mult_Buf[54].Weight_n = Wgt_6_250;
         Mult_Buf[55].Feature_n = FeatureBuf_251;
         Mult_Buf[55].Weight_n = Wgt_6_251;
         Mult_Buf[56].Feature_n = FeatureBuf_252;
         Mult_Buf[56].Weight_n = Wgt_6_252;
         Mult_Buf[57].Feature_n = FeatureBuf_253;
         Mult_Buf[57].Weight_n = Wgt_6_253;
         Mult_Buf[58].Feature_n = FeatureBuf_254;
         Mult_Buf[58].Weight_n = Wgt_6_254;
         Mult_Buf[59].Feature_n = FeatureBuf_255;
         Mult_Buf[59].Weight_n = Wgt_6_255;
         Mult_Buf[60].Feature_n = FeatureBuf_256;
         Mult_Buf[60].Weight_n = Wgt_6_256;
         Mult_Buf[61].Feature_n = FeatureBuf_257;
         Mult_Buf[61].Weight_n = Wgt_6_257;
         Mult_Buf[62].Feature_n = FeatureBuf_258;
         Mult_Buf[62].Weight_n = Wgt_6_258;
         Mult_Buf[63].Feature_n = FeatureBuf_259;
         Mult_Buf[63].Weight_n = Wgt_6_259;
         Mult_Buf[64].Feature_n = FeatureBuf_260;
         Mult_Buf[64].Weight_n = Wgt_6_260;
         Mult_Buf[65].Feature_n = FeatureBuf_261;
         Mult_Buf[65].Weight_n = Wgt_6_261;
         Mult_Buf[66].Feature_n = FeatureBuf_262;
         Mult_Buf[66].Weight_n = Wgt_6_262;
         Mult_Buf[67].Feature_n = FeatureBuf_263;
         Mult_Buf[67].Weight_n = Wgt_6_263;
         Mult_Buf[68].Feature_n = FeatureBuf_264;
         Mult_Buf[68].Weight_n = Wgt_6_264;
         Mult_Buf[69].Feature_n = FeatureBuf_265;
         Mult_Buf[69].Weight_n = Wgt_6_265;
         Mult_Buf[70].Feature_n = FeatureBuf_266;
         Mult_Buf[70].Weight_n = Wgt_6_266;
         Mult_Buf[71].Feature_n = FeatureBuf_267;
         Mult_Buf[71].Weight_n = Wgt_6_267;
         Mult_Buf[72].Feature_n = FeatureBuf_268;
         Mult_Buf[72].Weight_n = Wgt_6_268;
         Mult_Buf[73].Feature_n = FeatureBuf_269;
         Mult_Buf[73].Weight_n = Wgt_6_269;
         Mult_Buf[74].Feature_n = FeatureBuf_270;
         Mult_Buf[74].Weight_n = Wgt_6_270;
         Mult_Buf[75].Feature_n = FeatureBuf_271;
         Mult_Buf[75].Weight_n = Wgt_6_271;
         Mult_Buf[76].Feature_n = FeatureBuf_272;
         Mult_Buf[76].Weight_n = Wgt_6_272;
         Mult_Buf[77].Feature_n = FeatureBuf_273;
         Mult_Buf[77].Weight_n = Wgt_6_273;
         Mult_Buf[78].Feature_n = FeatureBuf_274;
         Mult_Buf[78].Weight_n = Wgt_6_274;
         Mult_Buf[79].Feature_n = FeatureBuf_275;
         Mult_Buf[79].Weight_n = Wgt_6_275;
         Mult_Buf[80].Feature_n = FeatureBuf_276;
         Mult_Buf[80].Weight_n = Wgt_6_276;
         Mult_Buf[81].Feature_n = FeatureBuf_277;
         Mult_Buf[81].Weight_n = Wgt_6_277;
         Mult_Buf[82].Feature_n = FeatureBuf_278;
         Mult_Buf[82].Weight_n = Wgt_6_278;
         Mult_Buf[83].Feature_n = FeatureBuf_279;
         Mult_Buf[83].Weight_n = Wgt_6_279;
         Mult_Buf[84].Feature_n = FeatureBuf_280;
         Mult_Buf[84].Weight_n = Wgt_6_280;
         Mult_Buf[85].Feature_n = FeatureBuf_281;
         Mult_Buf[85].Weight_n = Wgt_6_281;
         Mult_Buf[86].Feature_n = FeatureBuf_282;
         Mult_Buf[86].Weight_n = Wgt_6_282;
         Mult_Buf[87].Feature_n = FeatureBuf_283;
         Mult_Buf[87].Weight_n = Wgt_6_283;
         Mult_Buf[88].Feature_n = FeatureBuf_284;
         Mult_Buf[88].Weight_n = Wgt_6_284;
         Mult_Buf[89].Feature_n = FeatureBuf_285;
         Mult_Buf[89].Weight_n = Wgt_6_285;
         Mult_Buf[90].Feature_n = FeatureBuf_286;
         Mult_Buf[90].Weight_n = Wgt_6_286;
         Mult_Buf[91].Feature_n = FeatureBuf_287;
         Mult_Buf[91].Weight_n = Wgt_6_287;
         Mult_Buf[92].Feature_n = FeatureBuf_288;
         Mult_Buf[92].Weight_n = Wgt_6_288;
         Mult_Buf[93].Feature_n = FeatureBuf_289;
         Mult_Buf[93].Weight_n = Wgt_6_289;
         Mult_Buf[94].Feature_n = FeatureBuf_290;
         Mult_Buf[94].Weight_n = Wgt_6_290;
         Mult_Buf[95].Feature_n = FeatureBuf_291;
         Mult_Buf[95].Weight_n = Wgt_6_291;
         Mult_Buf[96].Feature_n = FeatureBuf_292;
         Mult_Buf[96].Weight_n = Wgt_6_292;
         Mult_Buf[97].Feature_n = FeatureBuf_293;
         Mult_Buf[97].Weight_n = Wgt_6_293;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     //Collect Partial result form Adder
         Res_3_4_n = Part_Res;
     end
    53:begin
     nxt_state = 54;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_294;
         Mult_Buf[0].Weight_n = Wgt_6_294;
         Mult_Buf[1].Feature_n = FeatureBuf_295;
         Mult_Buf[1].Weight_n = Wgt_6_295;
         Mult_Buf[2].Feature_n = FeatureBuf_296;
         Mult_Buf[2].Weight_n = Wgt_6_296;
         Mult_Buf[3].Feature_n = FeatureBuf_297;
         Mult_Buf[3].Weight_n = Wgt_6_297;
         Mult_Buf[4].Feature_n = FeatureBuf_298;
         Mult_Buf[4].Weight_n = Wgt_6_298;
         Mult_Buf[5].Feature_n = FeatureBuf_299;
         Mult_Buf[5].Weight_n = Wgt_6_299;
         Mult_Buf[6].Feature_n = FeatureBuf_300;
         Mult_Buf[6].Weight_n = Wgt_6_300;
         Mult_Buf[7].Feature_n = FeatureBuf_301;
         Mult_Buf[7].Weight_n = Wgt_6_301;
         Mult_Buf[8].Feature_n = FeatureBuf_302;
         Mult_Buf[8].Weight_n = Wgt_6_302;
         Mult_Buf[9].Feature_n = FeatureBuf_303;
         Mult_Buf[9].Weight_n = Wgt_6_303;
         Mult_Buf[10].Feature_n = FeatureBuf_304;
         Mult_Buf[10].Weight_n = Wgt_6_304;
         Mult_Buf[11].Feature_n = FeatureBuf_305;
         Mult_Buf[11].Weight_n = Wgt_6_305;
         Mult_Buf[12].Feature_n = FeatureBuf_306;
         Mult_Buf[12].Weight_n = Wgt_6_306;
         Mult_Buf[13].Feature_n = FeatureBuf_307;
         Mult_Buf[13].Weight_n = Wgt_6_307;
         Mult_Buf[14].Feature_n = FeatureBuf_308;
         Mult_Buf[14].Weight_n = Wgt_6_308;
         Mult_Buf[15].Feature_n = FeatureBuf_309;
         Mult_Buf[15].Weight_n = Wgt_6_309;
         Mult_Buf[16].Feature_n = FeatureBuf_310;
         Mult_Buf[16].Weight_n = Wgt_6_310;
         Mult_Buf[17].Feature_n = FeatureBuf_311;
         Mult_Buf[17].Weight_n = Wgt_6_311;
         Mult_Buf[18].Feature_n = FeatureBuf_312;
         Mult_Buf[18].Weight_n = Wgt_6_312;
         Mult_Buf[19].Feature_n = FeatureBuf_313;
         Mult_Buf[19].Weight_n = Wgt_6_313;
         Mult_Buf[20].Feature_n = FeatureBuf_314;
         Mult_Buf[20].Weight_n = Wgt_6_314;
         Mult_Buf[21].Feature_n = FeatureBuf_315;
         Mult_Buf[21].Weight_n = Wgt_6_315;
         Mult_Buf[22].Feature_n = FeatureBuf_316;
         Mult_Buf[22].Weight_n = Wgt_6_316;
         Mult_Buf[23].Feature_n = FeatureBuf_317;
         Mult_Buf[23].Weight_n = Wgt_6_317;
         Mult_Buf[24].Feature_n = FeatureBuf_318;
         Mult_Buf[24].Weight_n = Wgt_6_318;
         Mult_Buf[25].Feature_n = FeatureBuf_319;
         Mult_Buf[25].Weight_n = Wgt_6_319;
         Mult_Buf[26].Feature_n = FeatureBuf_320;
         Mult_Buf[26].Weight_n = Wgt_6_320;
         Mult_Buf[27].Feature_n = FeatureBuf_321;
         Mult_Buf[27].Weight_n = Wgt_6_321;
         Mult_Buf[28].Feature_n = FeatureBuf_322;
         Mult_Buf[28].Weight_n = Wgt_6_322;
         Mult_Buf[29].Feature_n = FeatureBuf_323;
         Mult_Buf[29].Weight_n = Wgt_6_323;
         Mult_Buf[30].Feature_n = FeatureBuf_324;
         Mult_Buf[30].Weight_n = Wgt_6_324;
         Mult_Buf[31].Feature_n = FeatureBuf_325;
         Mult_Buf[31].Weight_n = Wgt_6_325;
         Mult_Buf[32].Feature_n = FeatureBuf_326;
         Mult_Buf[32].Weight_n = Wgt_6_326;
         Mult_Buf[33].Feature_n = FeatureBuf_327;
         Mult_Buf[33].Weight_n = Wgt_6_327;
         Mult_Buf[34].Feature_n = FeatureBuf_328;
         Mult_Buf[34].Weight_n = Wgt_6_328;
         Mult_Buf[35].Feature_n = FeatureBuf_329;
         Mult_Buf[35].Weight_n = Wgt_6_329;
         Mult_Buf[36].Feature_n = FeatureBuf_330;
         Mult_Buf[36].Weight_n = Wgt_6_330;
         Mult_Buf[37].Feature_n = FeatureBuf_331;
         Mult_Buf[37].Weight_n = Wgt_6_331;
         Mult_Buf[38].Feature_n = FeatureBuf_332;
         Mult_Buf[38].Weight_n = Wgt_6_332;
         Mult_Buf[39].Feature_n = FeatureBuf_333;
         Mult_Buf[39].Weight_n = Wgt_6_333;
         Mult_Buf[40].Feature_n = FeatureBuf_334;
         Mult_Buf[40].Weight_n = Wgt_6_334;
         Mult_Buf[41].Feature_n = FeatureBuf_335;
         Mult_Buf[41].Weight_n = Wgt_6_335;
         Mult_Buf[42].Feature_n = FeatureBuf_336;
         Mult_Buf[42].Weight_n = Wgt_6_336;
         Mult_Buf[43].Feature_n = FeatureBuf_337;
         Mult_Buf[43].Weight_n = Wgt_6_337;
         Mult_Buf[44].Feature_n = FeatureBuf_338;
         Mult_Buf[44].Weight_n = Wgt_6_338;
         Mult_Buf[45].Feature_n = FeatureBuf_339;
         Mult_Buf[45].Weight_n = Wgt_6_339;
         Mult_Buf[46].Feature_n = FeatureBuf_340;
         Mult_Buf[46].Weight_n = Wgt_6_340;
         Mult_Buf[47].Feature_n = FeatureBuf_341;
         Mult_Buf[47].Weight_n = Wgt_6_341;
         Mult_Buf[48].Feature_n = FeatureBuf_342;
         Mult_Buf[48].Weight_n = Wgt_6_342;
         Mult_Buf[49].Feature_n = FeatureBuf_343;
         Mult_Buf[49].Weight_n = Wgt_6_343;
         Mult_Buf[50].Feature_n = FeatureBuf_344;
         Mult_Buf[50].Weight_n = Wgt_6_344;
         Mult_Buf[51].Feature_n = FeatureBuf_345;
         Mult_Buf[51].Weight_n = Wgt_6_345;
         Mult_Buf[52].Feature_n = FeatureBuf_346;
         Mult_Buf[52].Weight_n = Wgt_6_346;
         Mult_Buf[53].Feature_n = FeatureBuf_347;
         Mult_Buf[53].Weight_n = Wgt_6_347;
         Mult_Buf[54].Feature_n = FeatureBuf_348;
         Mult_Buf[54].Weight_n = Wgt_6_348;
         Mult_Buf[55].Feature_n = FeatureBuf_349;
         Mult_Buf[55].Weight_n = Wgt_6_349;
         Mult_Buf[56].Feature_n = FeatureBuf_350;
         Mult_Buf[56].Weight_n = Wgt_6_350;
         Mult_Buf[57].Feature_n = FeatureBuf_351;
         Mult_Buf[57].Weight_n = Wgt_6_351;
         Mult_Buf[58].Feature_n = FeatureBuf_352;
         Mult_Buf[58].Weight_n = Wgt_6_352;
         Mult_Buf[59].Feature_n = FeatureBuf_353;
         Mult_Buf[59].Weight_n = Wgt_6_353;
         Mult_Buf[60].Feature_n = FeatureBuf_354;
         Mult_Buf[60].Weight_n = Wgt_6_354;
         Mult_Buf[61].Feature_n = FeatureBuf_355;
         Mult_Buf[61].Weight_n = Wgt_6_355;
         Mult_Buf[62].Feature_n = FeatureBuf_356;
         Mult_Buf[62].Weight_n = Wgt_6_356;
         Mult_Buf[63].Feature_n = FeatureBuf_357;
         Mult_Buf[63].Weight_n = Wgt_6_357;
         Mult_Buf[64].Feature_n = FeatureBuf_358;
         Mult_Buf[64].Weight_n = Wgt_6_358;
         Mult_Buf[65].Feature_n = FeatureBuf_359;
         Mult_Buf[65].Weight_n = Wgt_6_359;
         Mult_Buf[66].Feature_n = FeatureBuf_360;
         Mult_Buf[66].Weight_n = Wgt_6_360;
         Mult_Buf[67].Feature_n = FeatureBuf_361;
         Mult_Buf[67].Weight_n = Wgt_6_361;
         Mult_Buf[68].Feature_n = FeatureBuf_362;
         Mult_Buf[68].Weight_n = Wgt_6_362;
         Mult_Buf[69].Feature_n = FeatureBuf_363;
         Mult_Buf[69].Weight_n = Wgt_6_363;
         Mult_Buf[70].Feature_n = FeatureBuf_364;
         Mult_Buf[70].Weight_n = Wgt_6_364;
         Mult_Buf[71].Feature_n = FeatureBuf_365;
         Mult_Buf[71].Weight_n = Wgt_6_365;
         Mult_Buf[72].Feature_n = FeatureBuf_366;
         Mult_Buf[72].Weight_n = Wgt_6_366;
         Mult_Buf[73].Feature_n = FeatureBuf_367;
         Mult_Buf[73].Weight_n = Wgt_6_367;
         Mult_Buf[74].Feature_n = FeatureBuf_368;
         Mult_Buf[74].Weight_n = Wgt_6_368;
         Mult_Buf[75].Feature_n = FeatureBuf_369;
         Mult_Buf[75].Weight_n = Wgt_6_369;
         Mult_Buf[76].Feature_n = FeatureBuf_370;
         Mult_Buf[76].Weight_n = Wgt_6_370;
         Mult_Buf[77].Feature_n = FeatureBuf_371;
         Mult_Buf[77].Weight_n = Wgt_6_371;
         Mult_Buf[78].Feature_n = FeatureBuf_372;
         Mult_Buf[78].Weight_n = Wgt_6_372;
         Mult_Buf[79].Feature_n = FeatureBuf_373;
         Mult_Buf[79].Weight_n = Wgt_6_373;
         Mult_Buf[80].Feature_n = FeatureBuf_374;
         Mult_Buf[80].Weight_n = Wgt_6_374;
         Mult_Buf[81].Feature_n = FeatureBuf_375;
         Mult_Buf[81].Weight_n = Wgt_6_375;
         Mult_Buf[82].Feature_n = FeatureBuf_376;
         Mult_Buf[82].Weight_n = Wgt_6_376;
         Mult_Buf[83].Feature_n = FeatureBuf_377;
         Mult_Buf[83].Weight_n = Wgt_6_377;
         Mult_Buf[84].Feature_n = FeatureBuf_378;
         Mult_Buf[84].Weight_n = Wgt_6_378;
         Mult_Buf[85].Feature_n = FeatureBuf_379;
         Mult_Buf[85].Weight_n = Wgt_6_379;
         Mult_Buf[86].Feature_n = FeatureBuf_380;
         Mult_Buf[86].Weight_n = Wgt_6_380;
         Mult_Buf[87].Feature_n = FeatureBuf_381;
         Mult_Buf[87].Weight_n = Wgt_6_381;
         Mult_Buf[88].Feature_n = FeatureBuf_382;
         Mult_Buf[88].Weight_n = Wgt_6_382;
         Mult_Buf[89].Feature_n = FeatureBuf_383;
         Mult_Buf[89].Weight_n = Wgt_6_383;
         Mult_Buf[90].Feature_n = FeatureBuf_384;
         Mult_Buf[90].Weight_n = Wgt_6_384;
         Mult_Buf[91].Feature_n = FeatureBuf_385;
         Mult_Buf[91].Weight_n = Wgt_6_385;
         Mult_Buf[92].Feature_n = FeatureBuf_386;
         Mult_Buf[92].Weight_n = Wgt_6_386;
         Mult_Buf[93].Feature_n = FeatureBuf_387;
         Mult_Buf[93].Weight_n = Wgt_6_387;
         Mult_Buf[94].Feature_n = FeatureBuf_388;
         Mult_Buf[94].Weight_n = Wgt_6_388;
         Mult_Buf[95].Feature_n = FeatureBuf_389;
         Mult_Buf[95].Weight_n = Wgt_6_389;
         Mult_Buf[96].Feature_n = FeatureBuf_390;
         Mult_Buf[96].Weight_n = Wgt_6_390;
         Mult_Buf[97].Feature_n = FeatureBuf_391;
         Mult_Buf[97].Weight_n = Wgt_6_391;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     //Collect Partial result form Adder
         Res_3_5_n = Part_Res;
     //Collect result from final Adder
         Res2_n = Final_Res;
     end
    54:begin
     nxt_state = 55;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_392;
         Mult_Buf[0].Weight_n = Wgt_6_392;
         Mult_Buf[1].Feature_n = FeatureBuf_393;
         Mult_Buf[1].Weight_n = Wgt_6_393;
         Mult_Buf[2].Feature_n = FeatureBuf_394;
         Mult_Buf[2].Weight_n = Wgt_6_394;
         Mult_Buf[3].Feature_n = FeatureBuf_395;
         Mult_Buf[3].Weight_n = Wgt_6_395;
         Mult_Buf[4].Feature_n = FeatureBuf_396;
         Mult_Buf[4].Weight_n = Wgt_6_396;
         Mult_Buf[5].Feature_n = FeatureBuf_397;
         Mult_Buf[5].Weight_n = Wgt_6_397;
         Mult_Buf[6].Feature_n = FeatureBuf_398;
         Mult_Buf[6].Weight_n = Wgt_6_398;
         Mult_Buf[7].Feature_n = FeatureBuf_399;
         Mult_Buf[7].Weight_n = Wgt_6_399;
         Mult_Buf[8].Feature_n = FeatureBuf_400;
         Mult_Buf[8].Weight_n = Wgt_6_400;
         Mult_Buf[9].Feature_n = FeatureBuf_401;
         Mult_Buf[9].Weight_n = Wgt_6_401;
         Mult_Buf[10].Feature_n = FeatureBuf_402;
         Mult_Buf[10].Weight_n = Wgt_6_402;
         Mult_Buf[11].Feature_n = FeatureBuf_403;
         Mult_Buf[11].Weight_n = Wgt_6_403;
         Mult_Buf[12].Feature_n = FeatureBuf_404;
         Mult_Buf[12].Weight_n = Wgt_6_404;
         Mult_Buf[13].Feature_n = FeatureBuf_405;
         Mult_Buf[13].Weight_n = Wgt_6_405;
         Mult_Buf[14].Feature_n = FeatureBuf_406;
         Mult_Buf[14].Weight_n = Wgt_6_406;
         Mult_Buf[15].Feature_n = FeatureBuf_407;
         Mult_Buf[15].Weight_n = Wgt_6_407;
         Mult_Buf[16].Feature_n = FeatureBuf_408;
         Mult_Buf[16].Weight_n = Wgt_6_408;
         Mult_Buf[17].Feature_n = FeatureBuf_409;
         Mult_Buf[17].Weight_n = Wgt_6_409;
         Mult_Buf[18].Feature_n = FeatureBuf_410;
         Mult_Buf[18].Weight_n = Wgt_6_410;
         Mult_Buf[19].Feature_n = FeatureBuf_411;
         Mult_Buf[19].Weight_n = Wgt_6_411;
         Mult_Buf[20].Feature_n = FeatureBuf_412;
         Mult_Buf[20].Weight_n = Wgt_6_412;
         Mult_Buf[21].Feature_n = FeatureBuf_413;
         Mult_Buf[21].Weight_n = Wgt_6_413;
         Mult_Buf[22].Feature_n = FeatureBuf_414;
         Mult_Buf[22].Weight_n = Wgt_6_414;
         Mult_Buf[23].Feature_n = FeatureBuf_415;
         Mult_Buf[23].Weight_n = Wgt_6_415;
         Mult_Buf[24].Feature_n = FeatureBuf_416;
         Mult_Buf[24].Weight_n = Wgt_6_416;
         Mult_Buf[25].Feature_n = FeatureBuf_417;
         Mult_Buf[25].Weight_n = Wgt_6_417;
         Mult_Buf[26].Feature_n = FeatureBuf_418;
         Mult_Buf[26].Weight_n = Wgt_6_418;
         Mult_Buf[27].Feature_n = FeatureBuf_419;
         Mult_Buf[27].Weight_n = Wgt_6_419;
         Mult_Buf[28].Feature_n = FeatureBuf_420;
         Mult_Buf[28].Weight_n = Wgt_6_420;
         Mult_Buf[29].Feature_n = FeatureBuf_421;
         Mult_Buf[29].Weight_n = Wgt_6_421;
         Mult_Buf[30].Feature_n = FeatureBuf_422;
         Mult_Buf[30].Weight_n = Wgt_6_422;
         Mult_Buf[31].Feature_n = FeatureBuf_423;
         Mult_Buf[31].Weight_n = Wgt_6_423;
         Mult_Buf[32].Feature_n = FeatureBuf_424;
         Mult_Buf[32].Weight_n = Wgt_6_424;
         Mult_Buf[33].Feature_n = FeatureBuf_425;
         Mult_Buf[33].Weight_n = Wgt_6_425;
         Mult_Buf[34].Feature_n = FeatureBuf_426;
         Mult_Buf[34].Weight_n = Wgt_6_426;
         Mult_Buf[35].Feature_n = FeatureBuf_427;
         Mult_Buf[35].Weight_n = Wgt_6_427;
         Mult_Buf[36].Feature_n = FeatureBuf_428;
         Mult_Buf[36].Weight_n = Wgt_6_428;
         Mult_Buf[37].Feature_n = FeatureBuf_429;
         Mult_Buf[37].Weight_n = Wgt_6_429;
         Mult_Buf[38].Feature_n = FeatureBuf_430;
         Mult_Buf[38].Weight_n = Wgt_6_430;
         Mult_Buf[39].Feature_n = FeatureBuf_431;
         Mult_Buf[39].Weight_n = Wgt_6_431;
         Mult_Buf[40].Feature_n = FeatureBuf_432;
         Mult_Buf[40].Weight_n = Wgt_6_432;
         Mult_Buf[41].Feature_n = FeatureBuf_433;
         Mult_Buf[41].Weight_n = Wgt_6_433;
         Mult_Buf[42].Feature_n = FeatureBuf_434;
         Mult_Buf[42].Weight_n = Wgt_6_434;
         Mult_Buf[43].Feature_n = FeatureBuf_435;
         Mult_Buf[43].Weight_n = Wgt_6_435;
         Mult_Buf[44].Feature_n = FeatureBuf_436;
         Mult_Buf[44].Weight_n = Wgt_6_436;
         Mult_Buf[45].Feature_n = FeatureBuf_437;
         Mult_Buf[45].Weight_n = Wgt_6_437;
         Mult_Buf[46].Feature_n = FeatureBuf_438;
         Mult_Buf[46].Weight_n = Wgt_6_438;
         Mult_Buf[47].Feature_n = FeatureBuf_439;
         Mult_Buf[47].Weight_n = Wgt_6_439;
         Mult_Buf[48].Feature_n = FeatureBuf_440;
         Mult_Buf[48].Weight_n = Wgt_6_440;
         Mult_Buf[49].Feature_n = FeatureBuf_441;
         Mult_Buf[49].Weight_n = Wgt_6_441;
         Mult_Buf[50].Feature_n = FeatureBuf_442;
         Mult_Buf[50].Weight_n = Wgt_6_442;
         Mult_Buf[51].Feature_n = FeatureBuf_443;
         Mult_Buf[51].Weight_n = Wgt_6_443;
         Mult_Buf[52].Feature_n = FeatureBuf_444;
         Mult_Buf[52].Weight_n = Wgt_6_444;
         Mult_Buf[53].Feature_n = FeatureBuf_445;
         Mult_Buf[53].Weight_n = Wgt_6_445;
         Mult_Buf[54].Feature_n = FeatureBuf_446;
         Mult_Buf[54].Weight_n = Wgt_6_446;
         Mult_Buf[55].Feature_n = FeatureBuf_447;
         Mult_Buf[55].Weight_n = Wgt_6_447;
         Mult_Buf[56].Feature_n = FeatureBuf_448;
         Mult_Buf[56].Weight_n = Wgt_6_448;
         Mult_Buf[57].Feature_n = FeatureBuf_449;
         Mult_Buf[57].Weight_n = Wgt_6_449;
         Mult_Buf[58].Feature_n = FeatureBuf_450;
         Mult_Buf[58].Weight_n = Wgt_6_450;
         Mult_Buf[59].Feature_n = FeatureBuf_451;
         Mult_Buf[59].Weight_n = Wgt_6_451;
         Mult_Buf[60].Feature_n = FeatureBuf_452;
         Mult_Buf[60].Weight_n = Wgt_6_452;
         Mult_Buf[61].Feature_n = FeatureBuf_453;
         Mult_Buf[61].Weight_n = Wgt_6_453;
         Mult_Buf[62].Feature_n = FeatureBuf_454;
         Mult_Buf[62].Weight_n = Wgt_6_454;
         Mult_Buf[63].Feature_n = FeatureBuf_455;
         Mult_Buf[63].Weight_n = Wgt_6_455;
         Mult_Buf[64].Feature_n = FeatureBuf_456;
         Mult_Buf[64].Weight_n = Wgt_6_456;
         Mult_Buf[65].Feature_n = FeatureBuf_457;
         Mult_Buf[65].Weight_n = Wgt_6_457;
         Mult_Buf[66].Feature_n = FeatureBuf_458;
         Mult_Buf[66].Weight_n = Wgt_6_458;
         Mult_Buf[67].Feature_n = FeatureBuf_459;
         Mult_Buf[67].Weight_n = Wgt_6_459;
         Mult_Buf[68].Feature_n = FeatureBuf_460;
         Mult_Buf[68].Weight_n = Wgt_6_460;
         Mult_Buf[69].Feature_n = FeatureBuf_461;
         Mult_Buf[69].Weight_n = Wgt_6_461;
         Mult_Buf[70].Feature_n = FeatureBuf_462;
         Mult_Buf[70].Weight_n = Wgt_6_462;
         Mult_Buf[71].Feature_n = FeatureBuf_463;
         Mult_Buf[71].Weight_n = Wgt_6_463;
         Mult_Buf[72].Feature_n = FeatureBuf_464;
         Mult_Buf[72].Weight_n = Wgt_6_464;
         Mult_Buf[73].Feature_n = FeatureBuf_465;
         Mult_Buf[73].Weight_n = Wgt_6_465;
         Mult_Buf[74].Feature_n = FeatureBuf_466;
         Mult_Buf[74].Weight_n = Wgt_6_466;
         Mult_Buf[75].Feature_n = FeatureBuf_467;
         Mult_Buf[75].Weight_n = Wgt_6_467;
         Mult_Buf[76].Feature_n = FeatureBuf_468;
         Mult_Buf[76].Weight_n = Wgt_6_468;
         Mult_Buf[77].Feature_n = FeatureBuf_469;
         Mult_Buf[77].Weight_n = Wgt_6_469;
         Mult_Buf[78].Feature_n = FeatureBuf_470;
         Mult_Buf[78].Weight_n = Wgt_6_470;
         Mult_Buf[79].Feature_n = FeatureBuf_471;
         Mult_Buf[79].Weight_n = Wgt_6_471;
         Mult_Buf[80].Feature_n = FeatureBuf_472;
         Mult_Buf[80].Weight_n = Wgt_6_472;
         Mult_Buf[81].Feature_n = FeatureBuf_473;
         Mult_Buf[81].Weight_n = Wgt_6_473;
         Mult_Buf[82].Feature_n = FeatureBuf_474;
         Mult_Buf[82].Weight_n = Wgt_6_474;
         Mult_Buf[83].Feature_n = FeatureBuf_475;
         Mult_Buf[83].Weight_n = Wgt_6_475;
         Mult_Buf[84].Feature_n = FeatureBuf_476;
         Mult_Buf[84].Weight_n = Wgt_6_476;
         Mult_Buf[85].Feature_n = FeatureBuf_477;
         Mult_Buf[85].Weight_n = Wgt_6_477;
         Mult_Buf[86].Feature_n = FeatureBuf_478;
         Mult_Buf[86].Weight_n = Wgt_6_478;
         Mult_Buf[87].Feature_n = FeatureBuf_479;
         Mult_Buf[87].Weight_n = Wgt_6_479;
         Mult_Buf[88].Feature_n = FeatureBuf_480;
         Mult_Buf[88].Weight_n = Wgt_6_480;
         Mult_Buf[89].Feature_n = FeatureBuf_481;
         Mult_Buf[89].Weight_n = Wgt_6_481;
         Mult_Buf[90].Feature_n = FeatureBuf_482;
         Mult_Buf[90].Weight_n = Wgt_6_482;
         Mult_Buf[91].Feature_n = FeatureBuf_483;
         Mult_Buf[91].Weight_n = Wgt_6_483;
         Mult_Buf[92].Feature_n = FeatureBuf_484;
         Mult_Buf[92].Weight_n = Wgt_6_484;
         Mult_Buf[93].Feature_n = FeatureBuf_485;
         Mult_Buf[93].Weight_n = Wgt_6_485;
         Mult_Buf[94].Feature_n = FeatureBuf_486;
         Mult_Buf[94].Weight_n = Wgt_6_486;
         Mult_Buf[95].Feature_n = FeatureBuf_487;
         Mult_Buf[95].Weight_n = Wgt_6_487;
         Mult_Buf[96].Feature_n = FeatureBuf_488;
         Mult_Buf[96].Weight_n = Wgt_6_488;
         Mult_Buf[97].Feature_n = FeatureBuf_489;
         Mult_Buf[97].Weight_n = Wgt_6_489;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     //Collect Partial result form Adder
         Res_3_6_n = Part_Res;
     end
    55:begin
     nxt_state = 56;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_490;
         Mult_Buf[0].Weight_n = Wgt_6_490;
         Mult_Buf[1].Feature_n = FeatureBuf_491;
         Mult_Buf[1].Weight_n = Wgt_6_491;
         Mult_Buf[2].Feature_n = FeatureBuf_492;
         Mult_Buf[2].Weight_n = Wgt_6_492;
         Mult_Buf[3].Feature_n = FeatureBuf_493;
         Mult_Buf[3].Weight_n = Wgt_6_493;
         Mult_Buf[4].Feature_n = FeatureBuf_494;
         Mult_Buf[4].Weight_n = Wgt_6_494;
         Mult_Buf[5].Feature_n = FeatureBuf_495;
         Mult_Buf[5].Weight_n = Wgt_6_495;
         Mult_Buf[6].Feature_n = FeatureBuf_496;
         Mult_Buf[6].Weight_n = Wgt_6_496;
         Mult_Buf[7].Feature_n = FeatureBuf_497;
         Mult_Buf[7].Weight_n = Wgt_6_497;
         Mult_Buf[8].Feature_n = FeatureBuf_498;
         Mult_Buf[8].Weight_n = Wgt_6_498;
         Mult_Buf[9].Feature_n = FeatureBuf_499;
         Mult_Buf[9].Weight_n = Wgt_6_499;
         Mult_Buf[10].Feature_n = FeatureBuf_500;
         Mult_Buf[10].Weight_n = Wgt_6_500;
         Mult_Buf[11].Feature_n = FeatureBuf_501;
         Mult_Buf[11].Weight_n = Wgt_6_501;
         Mult_Buf[12].Feature_n = FeatureBuf_502;
         Mult_Buf[12].Weight_n = Wgt_6_502;
         Mult_Buf[13].Feature_n = FeatureBuf_503;
         Mult_Buf[13].Weight_n = Wgt_6_503;
         Mult_Buf[14].Feature_n = FeatureBuf_504;
         Mult_Buf[14].Weight_n = Wgt_6_504;
         Mult_Buf[15].Feature_n = FeatureBuf_505;
         Mult_Buf[15].Weight_n = Wgt_6_505;
         Mult_Buf[16].Feature_n = FeatureBuf_506;
         Mult_Buf[16].Weight_n = Wgt_6_506;
         Mult_Buf[17].Feature_n = FeatureBuf_507;
         Mult_Buf[17].Weight_n = Wgt_6_507;
         Mult_Buf[18].Feature_n = FeatureBuf_508;
         Mult_Buf[18].Weight_n = Wgt_6_508;
         Mult_Buf[19].Feature_n = FeatureBuf_509;
         Mult_Buf[19].Weight_n = Wgt_6_509;
         Mult_Buf[20].Feature_n = FeatureBuf_510;
         Mult_Buf[20].Weight_n = Wgt_6_510;
         Mult_Buf[21].Feature_n = FeatureBuf_511;
         Mult_Buf[21].Weight_n = Wgt_6_511;
         Mult_Buf[22].Feature_n = FeatureBuf_512;
         Mult_Buf[22].Weight_n = Wgt_6_512;
         Mult_Buf[23].Feature_n = FeatureBuf_513;
         Mult_Buf[23].Weight_n = Wgt_6_513;
         Mult_Buf[24].Feature_n = FeatureBuf_514;
         Mult_Buf[24].Weight_n = Wgt_6_514;
         Mult_Buf[25].Feature_n = FeatureBuf_515;
         Mult_Buf[25].Weight_n = Wgt_6_515;
         Mult_Buf[26].Feature_n = FeatureBuf_516;
         Mult_Buf[26].Weight_n = Wgt_6_516;
         Mult_Buf[27].Feature_n = FeatureBuf_517;
         Mult_Buf[27].Weight_n = Wgt_6_517;
         Mult_Buf[28].Feature_n = FeatureBuf_518;
         Mult_Buf[28].Weight_n = Wgt_6_518;
         Mult_Buf[29].Feature_n = FeatureBuf_519;
         Mult_Buf[29].Weight_n = Wgt_6_519;
         Mult_Buf[30].Feature_n = FeatureBuf_520;
         Mult_Buf[30].Weight_n = Wgt_6_520;
         Mult_Buf[31].Feature_n = FeatureBuf_521;
         Mult_Buf[31].Weight_n = Wgt_6_521;
         Mult_Buf[32].Feature_n = FeatureBuf_522;
         Mult_Buf[32].Weight_n = Wgt_6_522;
         Mult_Buf[33].Feature_n = FeatureBuf_523;
         Mult_Buf[33].Weight_n = Wgt_6_523;
         Mult_Buf[34].Feature_n = FeatureBuf_524;
         Mult_Buf[34].Weight_n = Wgt_6_524;
         Mult_Buf[35].Feature_n = FeatureBuf_525;
         Mult_Buf[35].Weight_n = Wgt_6_525;
         Mult_Buf[36].Feature_n = FeatureBuf_526;
         Mult_Buf[36].Weight_n = Wgt_6_526;
         Mult_Buf[37].Feature_n = FeatureBuf_527;
         Mult_Buf[37].Weight_n = Wgt_6_527;
         Mult_Buf[38].Feature_n = FeatureBuf_528;
         Mult_Buf[38].Weight_n = Wgt_6_528;
         Mult_Buf[39].Feature_n = FeatureBuf_529;
         Mult_Buf[39].Weight_n = Wgt_6_529;
         Mult_Buf[40].Feature_n = FeatureBuf_530;
         Mult_Buf[40].Weight_n = Wgt_6_530;
         Mult_Buf[41].Feature_n = FeatureBuf_531;
         Mult_Buf[41].Weight_n = Wgt_6_531;
         Mult_Buf[42].Feature_n = FeatureBuf_532;
         Mult_Buf[42].Weight_n = Wgt_6_532;
         Mult_Buf[43].Feature_n = FeatureBuf_533;
         Mult_Buf[43].Weight_n = Wgt_6_533;
         Mult_Buf[44].Feature_n = FeatureBuf_534;
         Mult_Buf[44].Weight_n = Wgt_6_534;
         Mult_Buf[45].Feature_n = FeatureBuf_535;
         Mult_Buf[45].Weight_n = Wgt_6_535;
         Mult_Buf[46].Feature_n = FeatureBuf_536;
         Mult_Buf[46].Weight_n = Wgt_6_536;
         Mult_Buf[47].Feature_n = FeatureBuf_537;
         Mult_Buf[47].Weight_n = Wgt_6_537;
         Mult_Buf[48].Feature_n = FeatureBuf_538;
         Mult_Buf[48].Weight_n = Wgt_6_538;
         Mult_Buf[49].Feature_n = FeatureBuf_539;
         Mult_Buf[49].Weight_n = Wgt_6_539;
         Mult_Buf[50].Feature_n = FeatureBuf_540;
         Mult_Buf[50].Weight_n = Wgt_6_540;
         Mult_Buf[51].Feature_n = FeatureBuf_541;
         Mult_Buf[51].Weight_n = Wgt_6_541;
         Mult_Buf[52].Feature_n = FeatureBuf_542;
         Mult_Buf[52].Weight_n = Wgt_6_542;
         Mult_Buf[53].Feature_n = FeatureBuf_543;
         Mult_Buf[53].Weight_n = Wgt_6_543;
         Mult_Buf[54].Feature_n = FeatureBuf_544;
         Mult_Buf[54].Weight_n = Wgt_6_544;
         Mult_Buf[55].Feature_n = FeatureBuf_545;
         Mult_Buf[55].Weight_n = Wgt_6_545;
         Mult_Buf[56].Feature_n = FeatureBuf_546;
         Mult_Buf[56].Weight_n = Wgt_6_546;
         Mult_Buf[57].Feature_n = FeatureBuf_547;
         Mult_Buf[57].Weight_n = Wgt_6_547;
         Mult_Buf[58].Feature_n = FeatureBuf_548;
         Mult_Buf[58].Weight_n = Wgt_6_548;
         Mult_Buf[59].Feature_n = FeatureBuf_549;
         Mult_Buf[59].Weight_n = Wgt_6_549;
         Mult_Buf[60].Feature_n = FeatureBuf_550;
         Mult_Buf[60].Weight_n = Wgt_6_550;
         Mult_Buf[61].Feature_n = FeatureBuf_551;
         Mult_Buf[61].Weight_n = Wgt_6_551;
         Mult_Buf[62].Feature_n = FeatureBuf_552;
         Mult_Buf[62].Weight_n = Wgt_6_552;
         Mult_Buf[63].Feature_n = FeatureBuf_553;
         Mult_Buf[63].Weight_n = Wgt_6_553;
         Mult_Buf[64].Feature_n = FeatureBuf_554;
         Mult_Buf[64].Weight_n = Wgt_6_554;
         Mult_Buf[65].Feature_n = FeatureBuf_555;
         Mult_Buf[65].Weight_n = Wgt_6_555;
         Mult_Buf[66].Feature_n = FeatureBuf_556;
         Mult_Buf[66].Weight_n = Wgt_6_556;
         Mult_Buf[67].Feature_n = FeatureBuf_557;
         Mult_Buf[67].Weight_n = Wgt_6_557;
         Mult_Buf[68].Feature_n = FeatureBuf_558;
         Mult_Buf[68].Weight_n = Wgt_6_558;
         Mult_Buf[69].Feature_n = FeatureBuf_559;
         Mult_Buf[69].Weight_n = Wgt_6_559;
         Mult_Buf[70].Feature_n = FeatureBuf_560;
         Mult_Buf[70].Weight_n = Wgt_6_560;
         Mult_Buf[71].Feature_n = FeatureBuf_561;
         Mult_Buf[71].Weight_n = Wgt_6_561;
         Mult_Buf[72].Feature_n = FeatureBuf_562;
         Mult_Buf[72].Weight_n = Wgt_6_562;
         Mult_Buf[73].Feature_n = FeatureBuf_563;
         Mult_Buf[73].Weight_n = Wgt_6_563;
         Mult_Buf[74].Feature_n = FeatureBuf_564;
         Mult_Buf[74].Weight_n = Wgt_6_564;
         Mult_Buf[75].Feature_n = FeatureBuf_565;
         Mult_Buf[75].Weight_n = Wgt_6_565;
         Mult_Buf[76].Feature_n = FeatureBuf_566;
         Mult_Buf[76].Weight_n = Wgt_6_566;
         Mult_Buf[77].Feature_n = FeatureBuf_567;
         Mult_Buf[77].Weight_n = Wgt_6_567;
         Mult_Buf[78].Feature_n = FeatureBuf_568;
         Mult_Buf[78].Weight_n = Wgt_6_568;
         Mult_Buf[79].Feature_n = FeatureBuf_569;
         Mult_Buf[79].Weight_n = Wgt_6_569;
         Mult_Buf[80].Feature_n = FeatureBuf_570;
         Mult_Buf[80].Weight_n = Wgt_6_570;
         Mult_Buf[81].Feature_n = FeatureBuf_571;
         Mult_Buf[81].Weight_n = Wgt_6_571;
         Mult_Buf[82].Feature_n = FeatureBuf_572;
         Mult_Buf[82].Weight_n = Wgt_6_572;
         Mult_Buf[83].Feature_n = FeatureBuf_573;
         Mult_Buf[83].Weight_n = Wgt_6_573;
         Mult_Buf[84].Feature_n = FeatureBuf_574;
         Mult_Buf[84].Weight_n = Wgt_6_574;
         Mult_Buf[85].Feature_n = FeatureBuf_575;
         Mult_Buf[85].Weight_n = Wgt_6_575;
         Mult_Buf[86].Feature_n = FeatureBuf_576;
         Mult_Buf[86].Weight_n = Wgt_6_576;
         Mult_Buf[87].Feature_n = FeatureBuf_577;
         Mult_Buf[87].Weight_n = Wgt_6_577;
         Mult_Buf[88].Feature_n = FeatureBuf_578;
         Mult_Buf[88].Weight_n = Wgt_6_578;
         Mult_Buf[89].Feature_n = FeatureBuf_579;
         Mult_Buf[89].Weight_n = Wgt_6_579;
         Mult_Buf[90].Feature_n = FeatureBuf_580;
         Mult_Buf[90].Weight_n = Wgt_6_580;
         Mult_Buf[91].Feature_n = FeatureBuf_581;
         Mult_Buf[91].Weight_n = Wgt_6_581;
         Mult_Buf[92].Feature_n = FeatureBuf_582;
         Mult_Buf[92].Weight_n = Wgt_6_582;
         Mult_Buf[93].Feature_n = FeatureBuf_583;
         Mult_Buf[93].Weight_n = Wgt_6_583;
         Mult_Buf[94].Feature_n = FeatureBuf_584;
         Mult_Buf[94].Weight_n = Wgt_6_584;
         Mult_Buf[95].Feature_n = FeatureBuf_585;
         Mult_Buf[95].Weight_n = Wgt_6_585;
         Mult_Buf[96].Feature_n = FeatureBuf_586;
         Mult_Buf[96].Weight_n = Wgt_6_586;
         Mult_Buf[97].Feature_n = FeatureBuf_587;
         Mult_Buf[97].Weight_n = Wgt_6_587;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     //Collect Partial result form Adder
         Res_3_7_n = Part_Res;
     //Feed to final Adder
         A1 = Part_Res;
         A2 = Res_3_6_n;
         A3 = Res_3_5_n;
         A4 = Res_3_4_n;
         A5 = Res_3_3_n;
         A6 = Res_3_2_n;
         A7 = Res_3_1_n;
         A8 = Res_3_0_n;
     end
    56:begin
     nxt_state = 57;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_588;
         Mult_Buf[0].Weight_n = Wgt_6_588;
         Mult_Buf[1].Feature_n = FeatureBuf_589;
         Mult_Buf[1].Weight_n = Wgt_6_589;
         Mult_Buf[2].Feature_n = FeatureBuf_590;
         Mult_Buf[2].Weight_n = Wgt_6_590;
         Mult_Buf[3].Feature_n = FeatureBuf_591;
         Mult_Buf[3].Weight_n = Wgt_6_591;
         Mult_Buf[4].Feature_n = FeatureBuf_592;
         Mult_Buf[4].Weight_n = Wgt_6_592;
         Mult_Buf[5].Feature_n = FeatureBuf_593;
         Mult_Buf[5].Weight_n = Wgt_6_593;
         Mult_Buf[6].Feature_n = FeatureBuf_594;
         Mult_Buf[6].Weight_n = Wgt_6_594;
         Mult_Buf[7].Feature_n = FeatureBuf_595;
         Mult_Buf[7].Weight_n = Wgt_6_595;
         Mult_Buf[8].Feature_n = FeatureBuf_596;
         Mult_Buf[8].Weight_n = Wgt_6_596;
         Mult_Buf[9].Feature_n = FeatureBuf_597;
         Mult_Buf[9].Weight_n = Wgt_6_597;
         Mult_Buf[10].Feature_n = FeatureBuf_598;
         Mult_Buf[10].Weight_n = Wgt_6_598;
         Mult_Buf[11].Feature_n = FeatureBuf_599;
         Mult_Buf[11].Weight_n = Wgt_6_599;
         Mult_Buf[12].Feature_n = FeatureBuf_600;
         Mult_Buf[12].Weight_n = Wgt_6_600;
         Mult_Buf[13].Feature_n = FeatureBuf_601;
         Mult_Buf[13].Weight_n = Wgt_6_601;
         Mult_Buf[14].Feature_n = FeatureBuf_602;
         Mult_Buf[14].Weight_n = Wgt_6_602;
         Mult_Buf[15].Feature_n = FeatureBuf_603;
         Mult_Buf[15].Weight_n = Wgt_6_603;
         Mult_Buf[16].Feature_n = FeatureBuf_604;
         Mult_Buf[16].Weight_n = Wgt_6_604;
         Mult_Buf[17].Feature_n = FeatureBuf_605;
         Mult_Buf[17].Weight_n = Wgt_6_605;
         Mult_Buf[18].Feature_n = FeatureBuf_606;
         Mult_Buf[18].Weight_n = Wgt_6_606;
         Mult_Buf[19].Feature_n = FeatureBuf_607;
         Mult_Buf[19].Weight_n = Wgt_6_607;
         Mult_Buf[20].Feature_n = FeatureBuf_608;
         Mult_Buf[20].Weight_n = Wgt_6_608;
         Mult_Buf[21].Feature_n = FeatureBuf_609;
         Mult_Buf[21].Weight_n = Wgt_6_609;
         Mult_Buf[22].Feature_n = FeatureBuf_610;
         Mult_Buf[22].Weight_n = Wgt_6_610;
         Mult_Buf[23].Feature_n = FeatureBuf_611;
         Mult_Buf[23].Weight_n = Wgt_6_611;
         Mult_Buf[24].Feature_n = FeatureBuf_612;
         Mult_Buf[24].Weight_n = Wgt_6_612;
         Mult_Buf[25].Feature_n = FeatureBuf_613;
         Mult_Buf[25].Weight_n = Wgt_6_613;
         Mult_Buf[26].Feature_n = FeatureBuf_614;
         Mult_Buf[26].Weight_n = Wgt_6_614;
         Mult_Buf[27].Feature_n = FeatureBuf_615;
         Mult_Buf[27].Weight_n = Wgt_6_615;
         Mult_Buf[28].Feature_n = FeatureBuf_616;
         Mult_Buf[28].Weight_n = Wgt_6_616;
         Mult_Buf[29].Feature_n = FeatureBuf_617;
         Mult_Buf[29].Weight_n = Wgt_6_617;
         Mult_Buf[30].Feature_n = FeatureBuf_618;
         Mult_Buf[30].Weight_n = Wgt_6_618;
         Mult_Buf[31].Feature_n = FeatureBuf_619;
         Mult_Buf[31].Weight_n = Wgt_6_619;
         Mult_Buf[32].Feature_n = FeatureBuf_620;
         Mult_Buf[32].Weight_n = Wgt_6_620;
         Mult_Buf[33].Feature_n = FeatureBuf_621;
         Mult_Buf[33].Weight_n = Wgt_6_621;
         Mult_Buf[34].Feature_n = FeatureBuf_622;
         Mult_Buf[34].Weight_n = Wgt_6_622;
         Mult_Buf[35].Feature_n = FeatureBuf_623;
         Mult_Buf[35].Weight_n = Wgt_6_623;
         Mult_Buf[36].Feature_n = FeatureBuf_624;
         Mult_Buf[36].Weight_n = Wgt_6_624;
         Mult_Buf[37].Feature_n = FeatureBuf_625;
         Mult_Buf[37].Weight_n = Wgt_6_625;
         Mult_Buf[38].Feature_n = FeatureBuf_626;
         Mult_Buf[38].Weight_n = Wgt_6_626;
         Mult_Buf[39].Feature_n = FeatureBuf_627;
         Mult_Buf[39].Weight_n = Wgt_6_627;
         Mult_Buf[40].Feature_n = FeatureBuf_628;
         Mult_Buf[40].Weight_n = Wgt_6_628;
         Mult_Buf[41].Feature_n = FeatureBuf_629;
         Mult_Buf[41].Weight_n = Wgt_6_629;
         Mult_Buf[42].Feature_n = FeatureBuf_630;
         Mult_Buf[42].Weight_n = Wgt_6_630;
         Mult_Buf[43].Feature_n = FeatureBuf_631;
         Mult_Buf[43].Weight_n = Wgt_6_631;
         Mult_Buf[44].Feature_n = FeatureBuf_632;
         Mult_Buf[44].Weight_n = Wgt_6_632;
         Mult_Buf[45].Feature_n = FeatureBuf_633;
         Mult_Buf[45].Weight_n = Wgt_6_633;
         Mult_Buf[46].Feature_n = FeatureBuf_634;
         Mult_Buf[46].Weight_n = Wgt_6_634;
         Mult_Buf[47].Feature_n = FeatureBuf_635;
         Mult_Buf[47].Weight_n = Wgt_6_635;
         Mult_Buf[48].Feature_n = FeatureBuf_636;
         Mult_Buf[48].Weight_n = Wgt_6_636;
         Mult_Buf[49].Feature_n = FeatureBuf_637;
         Mult_Buf[49].Weight_n = Wgt_6_637;
         Mult_Buf[50].Feature_n = FeatureBuf_638;
         Mult_Buf[50].Weight_n = Wgt_6_638;
         Mult_Buf[51].Feature_n = FeatureBuf_639;
         Mult_Buf[51].Weight_n = Wgt_6_639;
         Mult_Buf[52].Feature_n = FeatureBuf_640;
         Mult_Buf[52].Weight_n = Wgt_6_640;
         Mult_Buf[53].Feature_n = FeatureBuf_641;
         Mult_Buf[53].Weight_n = Wgt_6_641;
         Mult_Buf[54].Feature_n = FeatureBuf_642;
         Mult_Buf[54].Weight_n = Wgt_6_642;
         Mult_Buf[55].Feature_n = FeatureBuf_643;
         Mult_Buf[55].Weight_n = Wgt_6_643;
         Mult_Buf[56].Feature_n = FeatureBuf_644;
         Mult_Buf[56].Weight_n = Wgt_6_644;
         Mult_Buf[57].Feature_n = FeatureBuf_645;
         Mult_Buf[57].Weight_n = Wgt_6_645;
         Mult_Buf[58].Feature_n = FeatureBuf_646;
         Mult_Buf[58].Weight_n = Wgt_6_646;
         Mult_Buf[59].Feature_n = FeatureBuf_647;
         Mult_Buf[59].Weight_n = Wgt_6_647;
         Mult_Buf[60].Feature_n = FeatureBuf_648;
         Mult_Buf[60].Weight_n = Wgt_6_648;
         Mult_Buf[61].Feature_n = FeatureBuf_649;
         Mult_Buf[61].Weight_n = Wgt_6_649;
         Mult_Buf[62].Feature_n = FeatureBuf_650;
         Mult_Buf[62].Weight_n = Wgt_6_650;
         Mult_Buf[63].Feature_n = FeatureBuf_651;
         Mult_Buf[63].Weight_n = Wgt_6_651;
         Mult_Buf[64].Feature_n = FeatureBuf_652;
         Mult_Buf[64].Weight_n = Wgt_6_652;
         Mult_Buf[65].Feature_n = FeatureBuf_653;
         Mult_Buf[65].Weight_n = Wgt_6_653;
         Mult_Buf[66].Feature_n = FeatureBuf_654;
         Mult_Buf[66].Weight_n = Wgt_6_654;
         Mult_Buf[67].Feature_n = FeatureBuf_655;
         Mult_Buf[67].Weight_n = Wgt_6_655;
         Mult_Buf[68].Feature_n = FeatureBuf_656;
         Mult_Buf[68].Weight_n = Wgt_6_656;
         Mult_Buf[69].Feature_n = FeatureBuf_657;
         Mult_Buf[69].Weight_n = Wgt_6_657;
         Mult_Buf[70].Feature_n = FeatureBuf_658;
         Mult_Buf[70].Weight_n = Wgt_6_658;
         Mult_Buf[71].Feature_n = FeatureBuf_659;
         Mult_Buf[71].Weight_n = Wgt_6_659;
         Mult_Buf[72].Feature_n = FeatureBuf_660;
         Mult_Buf[72].Weight_n = Wgt_6_660;
         Mult_Buf[73].Feature_n = FeatureBuf_661;
         Mult_Buf[73].Weight_n = Wgt_6_661;
         Mult_Buf[74].Feature_n = FeatureBuf_662;
         Mult_Buf[74].Weight_n = Wgt_6_662;
         Mult_Buf[75].Feature_n = FeatureBuf_663;
         Mult_Buf[75].Weight_n = Wgt_6_663;
         Mult_Buf[76].Feature_n = FeatureBuf_664;
         Mult_Buf[76].Weight_n = Wgt_6_664;
         Mult_Buf[77].Feature_n = FeatureBuf_665;
         Mult_Buf[77].Weight_n = Wgt_6_665;
         Mult_Buf[78].Feature_n = FeatureBuf_666;
         Mult_Buf[78].Weight_n = Wgt_6_666;
         Mult_Buf[79].Feature_n = FeatureBuf_667;
         Mult_Buf[79].Weight_n = Wgt_6_667;
         Mult_Buf[80].Feature_n = FeatureBuf_668;
         Mult_Buf[80].Weight_n = Wgt_6_668;
         Mult_Buf[81].Feature_n = FeatureBuf_669;
         Mult_Buf[81].Weight_n = Wgt_6_669;
         Mult_Buf[82].Feature_n = FeatureBuf_670;
         Mult_Buf[82].Weight_n = Wgt_6_670;
         Mult_Buf[83].Feature_n = FeatureBuf_671;
         Mult_Buf[83].Weight_n = Wgt_6_671;
         Mult_Buf[84].Feature_n = FeatureBuf_672;
         Mult_Buf[84].Weight_n = Wgt_6_672;
         Mult_Buf[85].Feature_n = FeatureBuf_673;
         Mult_Buf[85].Weight_n = Wgt_6_673;
         Mult_Buf[86].Feature_n = FeatureBuf_674;
         Mult_Buf[86].Weight_n = Wgt_6_674;
         Mult_Buf[87].Feature_n = FeatureBuf_675;
         Mult_Buf[87].Weight_n = Wgt_6_675;
         Mult_Buf[88].Feature_n = FeatureBuf_676;
         Mult_Buf[88].Weight_n = Wgt_6_676;
         Mult_Buf[89].Feature_n = FeatureBuf_677;
         Mult_Buf[89].Weight_n = Wgt_6_677;
         Mult_Buf[90].Feature_n = FeatureBuf_678;
         Mult_Buf[90].Weight_n = Wgt_6_678;
         Mult_Buf[91].Feature_n = FeatureBuf_679;
         Mult_Buf[91].Weight_n = Wgt_6_679;
         Mult_Buf[92].Feature_n = FeatureBuf_680;
         Mult_Buf[92].Weight_n = Wgt_6_680;
         Mult_Buf[93].Feature_n = FeatureBuf_681;
         Mult_Buf[93].Weight_n = Wgt_6_681;
         Mult_Buf[94].Feature_n = FeatureBuf_682;
         Mult_Buf[94].Weight_n = Wgt_6_682;
         Mult_Buf[95].Feature_n = FeatureBuf_683;
         Mult_Buf[95].Weight_n = Wgt_6_683;
         Mult_Buf[96].Feature_n = FeatureBuf_684;
         Mult_Buf[96].Weight_n = Wgt_6_684;
         Mult_Buf[97].Feature_n = FeatureBuf_685;
         Mult_Buf[97].Weight_n = Wgt_6_685;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     //Collect Partial result form Adder
         Res_4_0_n = Part_Res;
     end
    57:begin
     nxt_state = 58;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_686;
         Mult_Buf[0].Weight_n = Wgt_6_686;
         Mult_Buf[1].Feature_n = FeatureBuf_687;
         Mult_Buf[1].Weight_n = Wgt_6_687;
         Mult_Buf[2].Feature_n = FeatureBuf_688;
         Mult_Buf[2].Weight_n = Wgt_6_688;
         Mult_Buf[3].Feature_n = FeatureBuf_689;
         Mult_Buf[3].Weight_n = Wgt_6_689;
         Mult_Buf[4].Feature_n = FeatureBuf_690;
         Mult_Buf[4].Weight_n = Wgt_6_690;
         Mult_Buf[5].Feature_n = FeatureBuf_691;
         Mult_Buf[5].Weight_n = Wgt_6_691;
         Mult_Buf[6].Feature_n = FeatureBuf_692;
         Mult_Buf[6].Weight_n = Wgt_6_692;
         Mult_Buf[7].Feature_n = FeatureBuf_693;
         Mult_Buf[7].Weight_n = Wgt_6_693;
         Mult_Buf[8].Feature_n = FeatureBuf_694;
         Mult_Buf[8].Weight_n = Wgt_6_694;
         Mult_Buf[9].Feature_n = FeatureBuf_695;
         Mult_Buf[9].Weight_n = Wgt_6_695;
         Mult_Buf[10].Feature_n = FeatureBuf_696;
         Mult_Buf[10].Weight_n = Wgt_6_696;
         Mult_Buf[11].Feature_n = FeatureBuf_697;
         Mult_Buf[11].Weight_n = Wgt_6_697;
         Mult_Buf[12].Feature_n = FeatureBuf_698;
         Mult_Buf[12].Weight_n = Wgt_6_698;
         Mult_Buf[13].Feature_n = FeatureBuf_699;
         Mult_Buf[13].Weight_n = Wgt_6_699;
         Mult_Buf[14].Feature_n = FeatureBuf_700;
         Mult_Buf[14].Weight_n = Wgt_6_700;
         Mult_Buf[15].Feature_n = FeatureBuf_701;
         Mult_Buf[15].Weight_n = Wgt_6_701;
         Mult_Buf[16].Feature_n = FeatureBuf_702;
         Mult_Buf[16].Weight_n = Wgt_6_702;
         Mult_Buf[17].Feature_n = FeatureBuf_703;
         Mult_Buf[17].Weight_n = Wgt_6_703;
         Mult_Buf[18].Feature_n = FeatureBuf_704;
         Mult_Buf[18].Weight_n = Wgt_6_704;
         Mult_Buf[19].Feature_n = FeatureBuf_705;
         Mult_Buf[19].Weight_n = Wgt_6_705;
         Mult_Buf[20].Feature_n = FeatureBuf_706;
         Mult_Buf[20].Weight_n = Wgt_6_706;
         Mult_Buf[21].Feature_n = FeatureBuf_707;
         Mult_Buf[21].Weight_n = Wgt_6_707;
         Mult_Buf[22].Feature_n = FeatureBuf_708;
         Mult_Buf[22].Weight_n = Wgt_6_708;
         Mult_Buf[23].Feature_n = FeatureBuf_709;
         Mult_Buf[23].Weight_n = Wgt_6_709;
         Mult_Buf[24].Feature_n = FeatureBuf_710;
         Mult_Buf[24].Weight_n = Wgt_6_710;
         Mult_Buf[25].Feature_n = FeatureBuf_711;
         Mult_Buf[25].Weight_n = Wgt_6_711;
         Mult_Buf[26].Feature_n = FeatureBuf_712;
         Mult_Buf[26].Weight_n = Wgt_6_712;
         Mult_Buf[27].Feature_n = FeatureBuf_713;
         Mult_Buf[27].Weight_n = Wgt_6_713;
         Mult_Buf[28].Feature_n = FeatureBuf_714;
         Mult_Buf[28].Weight_n = Wgt_6_714;
         Mult_Buf[29].Feature_n = FeatureBuf_715;
         Mult_Buf[29].Weight_n = Wgt_6_715;
         Mult_Buf[30].Feature_n = FeatureBuf_716;
         Mult_Buf[30].Weight_n = Wgt_6_716;
         Mult_Buf[31].Feature_n = FeatureBuf_717;
         Mult_Buf[31].Weight_n = Wgt_6_717;
         Mult_Buf[32].Feature_n = FeatureBuf_718;
         Mult_Buf[32].Weight_n = Wgt_6_718;
         Mult_Buf[33].Feature_n = FeatureBuf_719;
         Mult_Buf[33].Weight_n = Wgt_6_719;
         Mult_Buf[34].Feature_n = FeatureBuf_720;
         Mult_Buf[34].Weight_n = Wgt_6_720;
         Mult_Buf[35].Feature_n = FeatureBuf_721;
         Mult_Buf[35].Weight_n = Wgt_6_721;
         Mult_Buf[36].Feature_n = FeatureBuf_722;
         Mult_Buf[36].Weight_n = Wgt_6_722;
         Mult_Buf[37].Feature_n = FeatureBuf_723;
         Mult_Buf[37].Weight_n = Wgt_6_723;
         Mult_Buf[38].Feature_n = FeatureBuf_724;
         Mult_Buf[38].Weight_n = Wgt_6_724;
         Mult_Buf[39].Feature_n = FeatureBuf_725;
         Mult_Buf[39].Weight_n = Wgt_6_725;
         Mult_Buf[40].Feature_n = FeatureBuf_726;
         Mult_Buf[40].Weight_n = Wgt_6_726;
         Mult_Buf[41].Feature_n = FeatureBuf_727;
         Mult_Buf[41].Weight_n = Wgt_6_727;
         Mult_Buf[42].Feature_n = FeatureBuf_728;
         Mult_Buf[42].Weight_n = Wgt_6_728;
         Mult_Buf[43].Feature_n = FeatureBuf_729;
         Mult_Buf[43].Weight_n = Wgt_6_729;
         Mult_Buf[44].Feature_n = FeatureBuf_730;
         Mult_Buf[44].Weight_n = Wgt_6_730;
         Mult_Buf[45].Feature_n = FeatureBuf_731;
         Mult_Buf[45].Weight_n = Wgt_6_731;
         Mult_Buf[46].Feature_n = FeatureBuf_732;
         Mult_Buf[46].Weight_n = Wgt_6_732;
         Mult_Buf[47].Feature_n = FeatureBuf_733;
         Mult_Buf[47].Weight_n = Wgt_6_733;
         Mult_Buf[48].Feature_n = FeatureBuf_734;
         Mult_Buf[48].Weight_n = Wgt_6_734;
         Mult_Buf[49].Feature_n = FeatureBuf_735;
         Mult_Buf[49].Weight_n = Wgt_6_735;
         Mult_Buf[50].Feature_n = FeatureBuf_736;
         Mult_Buf[50].Weight_n = Wgt_6_736;
         Mult_Buf[51].Feature_n = FeatureBuf_737;
         Mult_Buf[51].Weight_n = Wgt_6_737;
         Mult_Buf[52].Feature_n = FeatureBuf_738;
         Mult_Buf[52].Weight_n = Wgt_6_738;
         Mult_Buf[53].Feature_n = FeatureBuf_739;
         Mult_Buf[53].Weight_n = Wgt_6_739;
         Mult_Buf[54].Feature_n = FeatureBuf_740;
         Mult_Buf[54].Weight_n = Wgt_6_740;
         Mult_Buf[55].Feature_n = FeatureBuf_741;
         Mult_Buf[55].Weight_n = Wgt_6_741;
         Mult_Buf[56].Feature_n = FeatureBuf_742;
         Mult_Buf[56].Weight_n = Wgt_6_742;
         Mult_Buf[57].Feature_n = FeatureBuf_743;
         Mult_Buf[57].Weight_n = Wgt_6_743;
         Mult_Buf[58].Feature_n = FeatureBuf_744;
         Mult_Buf[58].Weight_n = Wgt_6_744;
         Mult_Buf[59].Feature_n = FeatureBuf_745;
         Mult_Buf[59].Weight_n = Wgt_6_745;
         Mult_Buf[60].Feature_n = FeatureBuf_746;
         Mult_Buf[60].Weight_n = Wgt_6_746;
         Mult_Buf[61].Feature_n = FeatureBuf_747;
         Mult_Buf[61].Weight_n = Wgt_6_747;
         Mult_Buf[62].Feature_n = FeatureBuf_748;
         Mult_Buf[62].Weight_n = Wgt_6_748;
         Mult_Buf[63].Feature_n = FeatureBuf_749;
         Mult_Buf[63].Weight_n = Wgt_6_749;
         Mult_Buf[64].Feature_n = FeatureBuf_750;
         Mult_Buf[64].Weight_n = Wgt_6_750;
         Mult_Buf[65].Feature_n = FeatureBuf_751;
         Mult_Buf[65].Weight_n = Wgt_6_751;
         Mult_Buf[66].Feature_n = FeatureBuf_752;
         Mult_Buf[66].Weight_n = Wgt_6_752;
         Mult_Buf[67].Feature_n = FeatureBuf_753;
         Mult_Buf[67].Weight_n = Wgt_6_753;
         Mult_Buf[68].Feature_n = FeatureBuf_754;
         Mult_Buf[68].Weight_n = Wgt_6_754;
         Mult_Buf[69].Feature_n = FeatureBuf_755;
         Mult_Buf[69].Weight_n = Wgt_6_755;
         Mult_Buf[70].Feature_n = FeatureBuf_756;
         Mult_Buf[70].Weight_n = Wgt_6_756;
         Mult_Buf[71].Feature_n = FeatureBuf_757;
         Mult_Buf[71].Weight_n = Wgt_6_757;
         Mult_Buf[72].Feature_n = FeatureBuf_758;
         Mult_Buf[72].Weight_n = Wgt_6_758;
         Mult_Buf[73].Feature_n = FeatureBuf_759;
         Mult_Buf[73].Weight_n = Wgt_6_759;
         Mult_Buf[74].Feature_n = FeatureBuf_760;
         Mult_Buf[74].Weight_n = Wgt_6_760;
         Mult_Buf[75].Feature_n = FeatureBuf_761;
         Mult_Buf[75].Weight_n = Wgt_6_761;
         Mult_Buf[76].Feature_n = FeatureBuf_762;
         Mult_Buf[76].Weight_n = Wgt_6_762;
         Mult_Buf[77].Feature_n = FeatureBuf_763;
         Mult_Buf[77].Weight_n = Wgt_6_763;
         Mult_Buf[78].Feature_n = FeatureBuf_764;
         Mult_Buf[78].Weight_n = Wgt_6_764;
         Mult_Buf[79].Feature_n = FeatureBuf_765;
         Mult_Buf[79].Weight_n = Wgt_6_765;
         Mult_Buf[80].Feature_n = FeatureBuf_766;
         Mult_Buf[80].Weight_n = Wgt_6_766;
         Mult_Buf[81].Feature_n = FeatureBuf_767;
         Mult_Buf[81].Weight_n = Wgt_6_767;
         Mult_Buf[82].Feature_n = FeatureBuf_768;
         Mult_Buf[82].Weight_n = Wgt_6_768;
         Mult_Buf[83].Feature_n = FeatureBuf_769;
         Mult_Buf[83].Weight_n = Wgt_6_769;
         Mult_Buf[84].Feature_n = FeatureBuf_770;
         Mult_Buf[84].Weight_n = Wgt_6_770;
         Mult_Buf[85].Feature_n = FeatureBuf_771;
         Mult_Buf[85].Weight_n = Wgt_6_771;
         Mult_Buf[86].Feature_n = FeatureBuf_772;
         Mult_Buf[86].Weight_n = Wgt_6_772;
         Mult_Buf[87].Feature_n = FeatureBuf_773;
         Mult_Buf[87].Weight_n = Wgt_6_773;
         Mult_Buf[88].Feature_n = FeatureBuf_774;
         Mult_Buf[88].Weight_n = Wgt_6_774;
         Mult_Buf[89].Feature_n = FeatureBuf_775;
         Mult_Buf[89].Weight_n = Wgt_6_775;
         Mult_Buf[90].Feature_n = FeatureBuf_776;
         Mult_Buf[90].Weight_n = Wgt_6_776;
         Mult_Buf[91].Feature_n = FeatureBuf_777;
         Mult_Buf[91].Weight_n = Wgt_6_777;
         Mult_Buf[92].Feature_n = FeatureBuf_778;
         Mult_Buf[92].Weight_n = Wgt_6_778;
         Mult_Buf[93].Feature_n = FeatureBuf_779;
         Mult_Buf[93].Weight_n = Wgt_6_779;
         Mult_Buf[94].Feature_n = FeatureBuf_780;
         Mult_Buf[94].Weight_n = Wgt_6_780;
         Mult_Buf[95].Feature_n = FeatureBuf_781;
         Mult_Buf[95].Weight_n = Wgt_6_781;
         Mult_Buf[96].Feature_n = FeatureBuf_782;
         Mult_Buf[96].Weight_n = Wgt_6_782;
         Mult_Buf[97].Feature_n = FeatureBuf_783;
         Mult_Buf[97].Weight_n = Wgt_6_783;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     //Collect Partial result form Adder
         Res_4_1_n = Part_Res;
     end
    58:begin
     nxt_state = 59;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_0;
         Mult_Buf[0].Weight_n = Wgt_7_0;
         Mult_Buf[1].Feature_n = FeatureBuf_1;
         Mult_Buf[1].Weight_n = Wgt_7_1;
         Mult_Buf[2].Feature_n = FeatureBuf_2;
         Mult_Buf[2].Weight_n = Wgt_7_2;
         Mult_Buf[3].Feature_n = FeatureBuf_3;
         Mult_Buf[3].Weight_n = Wgt_7_3;
         Mult_Buf[4].Feature_n = FeatureBuf_4;
         Mult_Buf[4].Weight_n = Wgt_7_4;
         Mult_Buf[5].Feature_n = FeatureBuf_5;
         Mult_Buf[5].Weight_n = Wgt_7_5;
         Mult_Buf[6].Feature_n = FeatureBuf_6;
         Mult_Buf[6].Weight_n = Wgt_7_6;
         Mult_Buf[7].Feature_n = FeatureBuf_7;
         Mult_Buf[7].Weight_n = Wgt_7_7;
         Mult_Buf[8].Feature_n = FeatureBuf_8;
         Mult_Buf[8].Weight_n = Wgt_7_8;
         Mult_Buf[9].Feature_n = FeatureBuf_9;
         Mult_Buf[9].Weight_n = Wgt_7_9;
         Mult_Buf[10].Feature_n = FeatureBuf_10;
         Mult_Buf[10].Weight_n = Wgt_7_10;
         Mult_Buf[11].Feature_n = FeatureBuf_11;
         Mult_Buf[11].Weight_n = Wgt_7_11;
         Mult_Buf[12].Feature_n = FeatureBuf_12;
         Mult_Buf[12].Weight_n = Wgt_7_12;
         Mult_Buf[13].Feature_n = FeatureBuf_13;
         Mult_Buf[13].Weight_n = Wgt_7_13;
         Mult_Buf[14].Feature_n = FeatureBuf_14;
         Mult_Buf[14].Weight_n = Wgt_7_14;
         Mult_Buf[15].Feature_n = FeatureBuf_15;
         Mult_Buf[15].Weight_n = Wgt_7_15;
         Mult_Buf[16].Feature_n = FeatureBuf_16;
         Mult_Buf[16].Weight_n = Wgt_7_16;
         Mult_Buf[17].Feature_n = FeatureBuf_17;
         Mult_Buf[17].Weight_n = Wgt_7_17;
         Mult_Buf[18].Feature_n = FeatureBuf_18;
         Mult_Buf[18].Weight_n = Wgt_7_18;
         Mult_Buf[19].Feature_n = FeatureBuf_19;
         Mult_Buf[19].Weight_n = Wgt_7_19;
         Mult_Buf[20].Feature_n = FeatureBuf_20;
         Mult_Buf[20].Weight_n = Wgt_7_20;
         Mult_Buf[21].Feature_n = FeatureBuf_21;
         Mult_Buf[21].Weight_n = Wgt_7_21;
         Mult_Buf[22].Feature_n = FeatureBuf_22;
         Mult_Buf[22].Weight_n = Wgt_7_22;
         Mult_Buf[23].Feature_n = FeatureBuf_23;
         Mult_Buf[23].Weight_n = Wgt_7_23;
         Mult_Buf[24].Feature_n = FeatureBuf_24;
         Mult_Buf[24].Weight_n = Wgt_7_24;
         Mult_Buf[25].Feature_n = FeatureBuf_25;
         Mult_Buf[25].Weight_n = Wgt_7_25;
         Mult_Buf[26].Feature_n = FeatureBuf_26;
         Mult_Buf[26].Weight_n = Wgt_7_26;
         Mult_Buf[27].Feature_n = FeatureBuf_27;
         Mult_Buf[27].Weight_n = Wgt_7_27;
         Mult_Buf[28].Feature_n = FeatureBuf_28;
         Mult_Buf[28].Weight_n = Wgt_7_28;
         Mult_Buf[29].Feature_n = FeatureBuf_29;
         Mult_Buf[29].Weight_n = Wgt_7_29;
         Mult_Buf[30].Feature_n = FeatureBuf_30;
         Mult_Buf[30].Weight_n = Wgt_7_30;
         Mult_Buf[31].Feature_n = FeatureBuf_31;
         Mult_Buf[31].Weight_n = Wgt_7_31;
         Mult_Buf[32].Feature_n = FeatureBuf_32;
         Mult_Buf[32].Weight_n = Wgt_7_32;
         Mult_Buf[33].Feature_n = FeatureBuf_33;
         Mult_Buf[33].Weight_n = Wgt_7_33;
         Mult_Buf[34].Feature_n = FeatureBuf_34;
         Mult_Buf[34].Weight_n = Wgt_7_34;
         Mult_Buf[35].Feature_n = FeatureBuf_35;
         Mult_Buf[35].Weight_n = Wgt_7_35;
         Mult_Buf[36].Feature_n = FeatureBuf_36;
         Mult_Buf[36].Weight_n = Wgt_7_36;
         Mult_Buf[37].Feature_n = FeatureBuf_37;
         Mult_Buf[37].Weight_n = Wgt_7_37;
         Mult_Buf[38].Feature_n = FeatureBuf_38;
         Mult_Buf[38].Weight_n = Wgt_7_38;
         Mult_Buf[39].Feature_n = FeatureBuf_39;
         Mult_Buf[39].Weight_n = Wgt_7_39;
         Mult_Buf[40].Feature_n = FeatureBuf_40;
         Mult_Buf[40].Weight_n = Wgt_7_40;
         Mult_Buf[41].Feature_n = FeatureBuf_41;
         Mult_Buf[41].Weight_n = Wgt_7_41;
         Mult_Buf[42].Feature_n = FeatureBuf_42;
         Mult_Buf[42].Weight_n = Wgt_7_42;
         Mult_Buf[43].Feature_n = FeatureBuf_43;
         Mult_Buf[43].Weight_n = Wgt_7_43;
         Mult_Buf[44].Feature_n = FeatureBuf_44;
         Mult_Buf[44].Weight_n = Wgt_7_44;
         Mult_Buf[45].Feature_n = FeatureBuf_45;
         Mult_Buf[45].Weight_n = Wgt_7_45;
         Mult_Buf[46].Feature_n = FeatureBuf_46;
         Mult_Buf[46].Weight_n = Wgt_7_46;
         Mult_Buf[47].Feature_n = FeatureBuf_47;
         Mult_Buf[47].Weight_n = Wgt_7_47;
         Mult_Buf[48].Feature_n = FeatureBuf_48;
         Mult_Buf[48].Weight_n = Wgt_7_48;
         Mult_Buf[49].Feature_n = FeatureBuf_49;
         Mult_Buf[49].Weight_n = Wgt_7_49;
         Mult_Buf[50].Feature_n = FeatureBuf_50;
         Mult_Buf[50].Weight_n = Wgt_7_50;
         Mult_Buf[51].Feature_n = FeatureBuf_51;
         Mult_Buf[51].Weight_n = Wgt_7_51;
         Mult_Buf[52].Feature_n = FeatureBuf_52;
         Mult_Buf[52].Weight_n = Wgt_7_52;
         Mult_Buf[53].Feature_n = FeatureBuf_53;
         Mult_Buf[53].Weight_n = Wgt_7_53;
         Mult_Buf[54].Feature_n = FeatureBuf_54;
         Mult_Buf[54].Weight_n = Wgt_7_54;
         Mult_Buf[55].Feature_n = FeatureBuf_55;
         Mult_Buf[55].Weight_n = Wgt_7_55;
         Mult_Buf[56].Feature_n = FeatureBuf_56;
         Mult_Buf[56].Weight_n = Wgt_7_56;
         Mult_Buf[57].Feature_n = FeatureBuf_57;
         Mult_Buf[57].Weight_n = Wgt_7_57;
         Mult_Buf[58].Feature_n = FeatureBuf_58;
         Mult_Buf[58].Weight_n = Wgt_7_58;
         Mult_Buf[59].Feature_n = FeatureBuf_59;
         Mult_Buf[59].Weight_n = Wgt_7_59;
         Mult_Buf[60].Feature_n = FeatureBuf_60;
         Mult_Buf[60].Weight_n = Wgt_7_60;
         Mult_Buf[61].Feature_n = FeatureBuf_61;
         Mult_Buf[61].Weight_n = Wgt_7_61;
         Mult_Buf[62].Feature_n = FeatureBuf_62;
         Mult_Buf[62].Weight_n = Wgt_7_62;
         Mult_Buf[63].Feature_n = FeatureBuf_63;
         Mult_Buf[63].Weight_n = Wgt_7_63;
         Mult_Buf[64].Feature_n = FeatureBuf_64;
         Mult_Buf[64].Weight_n = Wgt_7_64;
         Mult_Buf[65].Feature_n = FeatureBuf_65;
         Mult_Buf[65].Weight_n = Wgt_7_65;
         Mult_Buf[66].Feature_n = FeatureBuf_66;
         Mult_Buf[66].Weight_n = Wgt_7_66;
         Mult_Buf[67].Feature_n = FeatureBuf_67;
         Mult_Buf[67].Weight_n = Wgt_7_67;
         Mult_Buf[68].Feature_n = FeatureBuf_68;
         Mult_Buf[68].Weight_n = Wgt_7_68;
         Mult_Buf[69].Feature_n = FeatureBuf_69;
         Mult_Buf[69].Weight_n = Wgt_7_69;
         Mult_Buf[70].Feature_n = FeatureBuf_70;
         Mult_Buf[70].Weight_n = Wgt_7_70;
         Mult_Buf[71].Feature_n = FeatureBuf_71;
         Mult_Buf[71].Weight_n = Wgt_7_71;
         Mult_Buf[72].Feature_n = FeatureBuf_72;
         Mult_Buf[72].Weight_n = Wgt_7_72;
         Mult_Buf[73].Feature_n = FeatureBuf_73;
         Mult_Buf[73].Weight_n = Wgt_7_73;
         Mult_Buf[74].Feature_n = FeatureBuf_74;
         Mult_Buf[74].Weight_n = Wgt_7_74;
         Mult_Buf[75].Feature_n = FeatureBuf_75;
         Mult_Buf[75].Weight_n = Wgt_7_75;
         Mult_Buf[76].Feature_n = FeatureBuf_76;
         Mult_Buf[76].Weight_n = Wgt_7_76;
         Mult_Buf[77].Feature_n = FeatureBuf_77;
         Mult_Buf[77].Weight_n = Wgt_7_77;
         Mult_Buf[78].Feature_n = FeatureBuf_78;
         Mult_Buf[78].Weight_n = Wgt_7_78;
         Mult_Buf[79].Feature_n = FeatureBuf_79;
         Mult_Buf[79].Weight_n = Wgt_7_79;
         Mult_Buf[80].Feature_n = FeatureBuf_80;
         Mult_Buf[80].Weight_n = Wgt_7_80;
         Mult_Buf[81].Feature_n = FeatureBuf_81;
         Mult_Buf[81].Weight_n = Wgt_7_81;
         Mult_Buf[82].Feature_n = FeatureBuf_82;
         Mult_Buf[82].Weight_n = Wgt_7_82;
         Mult_Buf[83].Feature_n = FeatureBuf_83;
         Mult_Buf[83].Weight_n = Wgt_7_83;
         Mult_Buf[84].Feature_n = FeatureBuf_84;
         Mult_Buf[84].Weight_n = Wgt_7_84;
         Mult_Buf[85].Feature_n = FeatureBuf_85;
         Mult_Buf[85].Weight_n = Wgt_7_85;
         Mult_Buf[86].Feature_n = FeatureBuf_86;
         Mult_Buf[86].Weight_n = Wgt_7_86;
         Mult_Buf[87].Feature_n = FeatureBuf_87;
         Mult_Buf[87].Weight_n = Wgt_7_87;
         Mult_Buf[88].Feature_n = FeatureBuf_88;
         Mult_Buf[88].Weight_n = Wgt_7_88;
         Mult_Buf[89].Feature_n = FeatureBuf_89;
         Mult_Buf[89].Weight_n = Wgt_7_89;
         Mult_Buf[90].Feature_n = FeatureBuf_90;
         Mult_Buf[90].Weight_n = Wgt_7_90;
         Mult_Buf[91].Feature_n = FeatureBuf_91;
         Mult_Buf[91].Weight_n = Wgt_7_91;
         Mult_Buf[92].Feature_n = FeatureBuf_92;
         Mult_Buf[92].Weight_n = Wgt_7_92;
         Mult_Buf[93].Feature_n = FeatureBuf_93;
         Mult_Buf[93].Weight_n = Wgt_7_93;
         Mult_Buf[94].Feature_n = FeatureBuf_94;
         Mult_Buf[94].Weight_n = Wgt_7_94;
         Mult_Buf[95].Feature_n = FeatureBuf_95;
         Mult_Buf[95].Weight_n = Wgt_7_95;
         Mult_Buf[96].Feature_n = FeatureBuf_96;
         Mult_Buf[96].Weight_n = Wgt_7_96;
         Mult_Buf[97].Feature_n = FeatureBuf_97;
         Mult_Buf[97].Weight_n = Wgt_7_97;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     //Collect Partial result form Adder
         Res_4_2_n = Part_Res;
     end
    59:begin
     nxt_state = 60;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_98;
         Mult_Buf[0].Weight_n = Wgt_7_98;
         Mult_Buf[1].Feature_n = FeatureBuf_99;
         Mult_Buf[1].Weight_n = Wgt_7_99;
         Mult_Buf[2].Feature_n = FeatureBuf_100;
         Mult_Buf[2].Weight_n = Wgt_7_100;
         Mult_Buf[3].Feature_n = FeatureBuf_101;
         Mult_Buf[3].Weight_n = Wgt_7_101;
         Mult_Buf[4].Feature_n = FeatureBuf_102;
         Mult_Buf[4].Weight_n = Wgt_7_102;
         Mult_Buf[5].Feature_n = FeatureBuf_103;
         Mult_Buf[5].Weight_n = Wgt_7_103;
         Mult_Buf[6].Feature_n = FeatureBuf_104;
         Mult_Buf[6].Weight_n = Wgt_7_104;
         Mult_Buf[7].Feature_n = FeatureBuf_105;
         Mult_Buf[7].Weight_n = Wgt_7_105;
         Mult_Buf[8].Feature_n = FeatureBuf_106;
         Mult_Buf[8].Weight_n = Wgt_7_106;
         Mult_Buf[9].Feature_n = FeatureBuf_107;
         Mult_Buf[9].Weight_n = Wgt_7_107;
         Mult_Buf[10].Feature_n = FeatureBuf_108;
         Mult_Buf[10].Weight_n = Wgt_7_108;
         Mult_Buf[11].Feature_n = FeatureBuf_109;
         Mult_Buf[11].Weight_n = Wgt_7_109;
         Mult_Buf[12].Feature_n = FeatureBuf_110;
         Mult_Buf[12].Weight_n = Wgt_7_110;
         Mult_Buf[13].Feature_n = FeatureBuf_111;
         Mult_Buf[13].Weight_n = Wgt_7_111;
         Mult_Buf[14].Feature_n = FeatureBuf_112;
         Mult_Buf[14].Weight_n = Wgt_7_112;
         Mult_Buf[15].Feature_n = FeatureBuf_113;
         Mult_Buf[15].Weight_n = Wgt_7_113;
         Mult_Buf[16].Feature_n = FeatureBuf_114;
         Mult_Buf[16].Weight_n = Wgt_7_114;
         Mult_Buf[17].Feature_n = FeatureBuf_115;
         Mult_Buf[17].Weight_n = Wgt_7_115;
         Mult_Buf[18].Feature_n = FeatureBuf_116;
         Mult_Buf[18].Weight_n = Wgt_7_116;
         Mult_Buf[19].Feature_n = FeatureBuf_117;
         Mult_Buf[19].Weight_n = Wgt_7_117;
         Mult_Buf[20].Feature_n = FeatureBuf_118;
         Mult_Buf[20].Weight_n = Wgt_7_118;
         Mult_Buf[21].Feature_n = FeatureBuf_119;
         Mult_Buf[21].Weight_n = Wgt_7_119;
         Mult_Buf[22].Feature_n = FeatureBuf_120;
         Mult_Buf[22].Weight_n = Wgt_7_120;
         Mult_Buf[23].Feature_n = FeatureBuf_121;
         Mult_Buf[23].Weight_n = Wgt_7_121;
         Mult_Buf[24].Feature_n = FeatureBuf_122;
         Mult_Buf[24].Weight_n = Wgt_7_122;
         Mult_Buf[25].Feature_n = FeatureBuf_123;
         Mult_Buf[25].Weight_n = Wgt_7_123;
         Mult_Buf[26].Feature_n = FeatureBuf_124;
         Mult_Buf[26].Weight_n = Wgt_7_124;
         Mult_Buf[27].Feature_n = FeatureBuf_125;
         Mult_Buf[27].Weight_n = Wgt_7_125;
         Mult_Buf[28].Feature_n = FeatureBuf_126;
         Mult_Buf[28].Weight_n = Wgt_7_126;
         Mult_Buf[29].Feature_n = FeatureBuf_127;
         Mult_Buf[29].Weight_n = Wgt_7_127;
         Mult_Buf[30].Feature_n = FeatureBuf_128;
         Mult_Buf[30].Weight_n = Wgt_7_128;
         Mult_Buf[31].Feature_n = FeatureBuf_129;
         Mult_Buf[31].Weight_n = Wgt_7_129;
         Mult_Buf[32].Feature_n = FeatureBuf_130;
         Mult_Buf[32].Weight_n = Wgt_7_130;
         Mult_Buf[33].Feature_n = FeatureBuf_131;
         Mult_Buf[33].Weight_n = Wgt_7_131;
         Mult_Buf[34].Feature_n = FeatureBuf_132;
         Mult_Buf[34].Weight_n = Wgt_7_132;
         Mult_Buf[35].Feature_n = FeatureBuf_133;
         Mult_Buf[35].Weight_n = Wgt_7_133;
         Mult_Buf[36].Feature_n = FeatureBuf_134;
         Mult_Buf[36].Weight_n = Wgt_7_134;
         Mult_Buf[37].Feature_n = FeatureBuf_135;
         Mult_Buf[37].Weight_n = Wgt_7_135;
         Mult_Buf[38].Feature_n = FeatureBuf_136;
         Mult_Buf[38].Weight_n = Wgt_7_136;
         Mult_Buf[39].Feature_n = FeatureBuf_137;
         Mult_Buf[39].Weight_n = Wgt_7_137;
         Mult_Buf[40].Feature_n = FeatureBuf_138;
         Mult_Buf[40].Weight_n = Wgt_7_138;
         Mult_Buf[41].Feature_n = FeatureBuf_139;
         Mult_Buf[41].Weight_n = Wgt_7_139;
         Mult_Buf[42].Feature_n = FeatureBuf_140;
         Mult_Buf[42].Weight_n = Wgt_7_140;
         Mult_Buf[43].Feature_n = FeatureBuf_141;
         Mult_Buf[43].Weight_n = Wgt_7_141;
         Mult_Buf[44].Feature_n = FeatureBuf_142;
         Mult_Buf[44].Weight_n = Wgt_7_142;
         Mult_Buf[45].Feature_n = FeatureBuf_143;
         Mult_Buf[45].Weight_n = Wgt_7_143;
         Mult_Buf[46].Feature_n = FeatureBuf_144;
         Mult_Buf[46].Weight_n = Wgt_7_144;
         Mult_Buf[47].Feature_n = FeatureBuf_145;
         Mult_Buf[47].Weight_n = Wgt_7_145;
         Mult_Buf[48].Feature_n = FeatureBuf_146;
         Mult_Buf[48].Weight_n = Wgt_7_146;
         Mult_Buf[49].Feature_n = FeatureBuf_147;
         Mult_Buf[49].Weight_n = Wgt_7_147;
         Mult_Buf[50].Feature_n = FeatureBuf_148;
         Mult_Buf[50].Weight_n = Wgt_7_148;
         Mult_Buf[51].Feature_n = FeatureBuf_149;
         Mult_Buf[51].Weight_n = Wgt_7_149;
         Mult_Buf[52].Feature_n = FeatureBuf_150;
         Mult_Buf[52].Weight_n = Wgt_7_150;
         Mult_Buf[53].Feature_n = FeatureBuf_151;
         Mult_Buf[53].Weight_n = Wgt_7_151;
         Mult_Buf[54].Feature_n = FeatureBuf_152;
         Mult_Buf[54].Weight_n = Wgt_7_152;
         Mult_Buf[55].Feature_n = FeatureBuf_153;
         Mult_Buf[55].Weight_n = Wgt_7_153;
         Mult_Buf[56].Feature_n = FeatureBuf_154;
         Mult_Buf[56].Weight_n = Wgt_7_154;
         Mult_Buf[57].Feature_n = FeatureBuf_155;
         Mult_Buf[57].Weight_n = Wgt_7_155;
         Mult_Buf[58].Feature_n = FeatureBuf_156;
         Mult_Buf[58].Weight_n = Wgt_7_156;
         Mult_Buf[59].Feature_n = FeatureBuf_157;
         Mult_Buf[59].Weight_n = Wgt_7_157;
         Mult_Buf[60].Feature_n = FeatureBuf_158;
         Mult_Buf[60].Weight_n = Wgt_7_158;
         Mult_Buf[61].Feature_n = FeatureBuf_159;
         Mult_Buf[61].Weight_n = Wgt_7_159;
         Mult_Buf[62].Feature_n = FeatureBuf_160;
         Mult_Buf[62].Weight_n = Wgt_7_160;
         Mult_Buf[63].Feature_n = FeatureBuf_161;
         Mult_Buf[63].Weight_n = Wgt_7_161;
         Mult_Buf[64].Feature_n = FeatureBuf_162;
         Mult_Buf[64].Weight_n = Wgt_7_162;
         Mult_Buf[65].Feature_n = FeatureBuf_163;
         Mult_Buf[65].Weight_n = Wgt_7_163;
         Mult_Buf[66].Feature_n = FeatureBuf_164;
         Mult_Buf[66].Weight_n = Wgt_7_164;
         Mult_Buf[67].Feature_n = FeatureBuf_165;
         Mult_Buf[67].Weight_n = Wgt_7_165;
         Mult_Buf[68].Feature_n = FeatureBuf_166;
         Mult_Buf[68].Weight_n = Wgt_7_166;
         Mult_Buf[69].Feature_n = FeatureBuf_167;
         Mult_Buf[69].Weight_n = Wgt_7_167;
         Mult_Buf[70].Feature_n = FeatureBuf_168;
         Mult_Buf[70].Weight_n = Wgt_7_168;
         Mult_Buf[71].Feature_n = FeatureBuf_169;
         Mult_Buf[71].Weight_n = Wgt_7_169;
         Mult_Buf[72].Feature_n = FeatureBuf_170;
         Mult_Buf[72].Weight_n = Wgt_7_170;
         Mult_Buf[73].Feature_n = FeatureBuf_171;
         Mult_Buf[73].Weight_n = Wgt_7_171;
         Mult_Buf[74].Feature_n = FeatureBuf_172;
         Mult_Buf[74].Weight_n = Wgt_7_172;
         Mult_Buf[75].Feature_n = FeatureBuf_173;
         Mult_Buf[75].Weight_n = Wgt_7_173;
         Mult_Buf[76].Feature_n = FeatureBuf_174;
         Mult_Buf[76].Weight_n = Wgt_7_174;
         Mult_Buf[77].Feature_n = FeatureBuf_175;
         Mult_Buf[77].Weight_n = Wgt_7_175;
         Mult_Buf[78].Feature_n = FeatureBuf_176;
         Mult_Buf[78].Weight_n = Wgt_7_176;
         Mult_Buf[79].Feature_n = FeatureBuf_177;
         Mult_Buf[79].Weight_n = Wgt_7_177;
         Mult_Buf[80].Feature_n = FeatureBuf_178;
         Mult_Buf[80].Weight_n = Wgt_7_178;
         Mult_Buf[81].Feature_n = FeatureBuf_179;
         Mult_Buf[81].Weight_n = Wgt_7_179;
         Mult_Buf[82].Feature_n = FeatureBuf_180;
         Mult_Buf[82].Weight_n = Wgt_7_180;
         Mult_Buf[83].Feature_n = FeatureBuf_181;
         Mult_Buf[83].Weight_n = Wgt_7_181;
         Mult_Buf[84].Feature_n = FeatureBuf_182;
         Mult_Buf[84].Weight_n = Wgt_7_182;
         Mult_Buf[85].Feature_n = FeatureBuf_183;
         Mult_Buf[85].Weight_n = Wgt_7_183;
         Mult_Buf[86].Feature_n = FeatureBuf_184;
         Mult_Buf[86].Weight_n = Wgt_7_184;
         Mult_Buf[87].Feature_n = FeatureBuf_185;
         Mult_Buf[87].Weight_n = Wgt_7_185;
         Mult_Buf[88].Feature_n = FeatureBuf_186;
         Mult_Buf[88].Weight_n = Wgt_7_186;
         Mult_Buf[89].Feature_n = FeatureBuf_187;
         Mult_Buf[89].Weight_n = Wgt_7_187;
         Mult_Buf[90].Feature_n = FeatureBuf_188;
         Mult_Buf[90].Weight_n = Wgt_7_188;
         Mult_Buf[91].Feature_n = FeatureBuf_189;
         Mult_Buf[91].Weight_n = Wgt_7_189;
         Mult_Buf[92].Feature_n = FeatureBuf_190;
         Mult_Buf[92].Weight_n = Wgt_7_190;
         Mult_Buf[93].Feature_n = FeatureBuf_191;
         Mult_Buf[93].Weight_n = Wgt_7_191;
         Mult_Buf[94].Feature_n = FeatureBuf_192;
         Mult_Buf[94].Weight_n = Wgt_7_192;
         Mult_Buf[95].Feature_n = FeatureBuf_193;
         Mult_Buf[95].Weight_n = Wgt_7_193;
         Mult_Buf[96].Feature_n = FeatureBuf_194;
         Mult_Buf[96].Weight_n = Wgt_7_194;
         Mult_Buf[97].Feature_n = FeatureBuf_195;
         Mult_Buf[97].Weight_n = Wgt_7_195;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     //Collect Partial result form Adder
         Res_4_3_n = Part_Res;
     end
    60:begin
     nxt_state = 61;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_196;
         Mult_Buf[0].Weight_n = Wgt_7_196;
         Mult_Buf[1].Feature_n = FeatureBuf_197;
         Mult_Buf[1].Weight_n = Wgt_7_197;
         Mult_Buf[2].Feature_n = FeatureBuf_198;
         Mult_Buf[2].Weight_n = Wgt_7_198;
         Mult_Buf[3].Feature_n = FeatureBuf_199;
         Mult_Buf[3].Weight_n = Wgt_7_199;
         Mult_Buf[4].Feature_n = FeatureBuf_200;
         Mult_Buf[4].Weight_n = Wgt_7_200;
         Mult_Buf[5].Feature_n = FeatureBuf_201;
         Mult_Buf[5].Weight_n = Wgt_7_201;
         Mult_Buf[6].Feature_n = FeatureBuf_202;
         Mult_Buf[6].Weight_n = Wgt_7_202;
         Mult_Buf[7].Feature_n = FeatureBuf_203;
         Mult_Buf[7].Weight_n = Wgt_7_203;
         Mult_Buf[8].Feature_n = FeatureBuf_204;
         Mult_Buf[8].Weight_n = Wgt_7_204;
         Mult_Buf[9].Feature_n = FeatureBuf_205;
         Mult_Buf[9].Weight_n = Wgt_7_205;
         Mult_Buf[10].Feature_n = FeatureBuf_206;
         Mult_Buf[10].Weight_n = Wgt_7_206;
         Mult_Buf[11].Feature_n = FeatureBuf_207;
         Mult_Buf[11].Weight_n = Wgt_7_207;
         Mult_Buf[12].Feature_n = FeatureBuf_208;
         Mult_Buf[12].Weight_n = Wgt_7_208;
         Mult_Buf[13].Feature_n = FeatureBuf_209;
         Mult_Buf[13].Weight_n = Wgt_7_209;
         Mult_Buf[14].Feature_n = FeatureBuf_210;
         Mult_Buf[14].Weight_n = Wgt_7_210;
         Mult_Buf[15].Feature_n = FeatureBuf_211;
         Mult_Buf[15].Weight_n = Wgt_7_211;
         Mult_Buf[16].Feature_n = FeatureBuf_212;
         Mult_Buf[16].Weight_n = Wgt_7_212;
         Mult_Buf[17].Feature_n = FeatureBuf_213;
         Mult_Buf[17].Weight_n = Wgt_7_213;
         Mult_Buf[18].Feature_n = FeatureBuf_214;
         Mult_Buf[18].Weight_n = Wgt_7_214;
         Mult_Buf[19].Feature_n = FeatureBuf_215;
         Mult_Buf[19].Weight_n = Wgt_7_215;
         Mult_Buf[20].Feature_n = FeatureBuf_216;
         Mult_Buf[20].Weight_n = Wgt_7_216;
         Mult_Buf[21].Feature_n = FeatureBuf_217;
         Mult_Buf[21].Weight_n = Wgt_7_217;
         Mult_Buf[22].Feature_n = FeatureBuf_218;
         Mult_Buf[22].Weight_n = Wgt_7_218;
         Mult_Buf[23].Feature_n = FeatureBuf_219;
         Mult_Buf[23].Weight_n = Wgt_7_219;
         Mult_Buf[24].Feature_n = FeatureBuf_220;
         Mult_Buf[24].Weight_n = Wgt_7_220;
         Mult_Buf[25].Feature_n = FeatureBuf_221;
         Mult_Buf[25].Weight_n = Wgt_7_221;
         Mult_Buf[26].Feature_n = FeatureBuf_222;
         Mult_Buf[26].Weight_n = Wgt_7_222;
         Mult_Buf[27].Feature_n = FeatureBuf_223;
         Mult_Buf[27].Weight_n = Wgt_7_223;
         Mult_Buf[28].Feature_n = FeatureBuf_224;
         Mult_Buf[28].Weight_n = Wgt_7_224;
         Mult_Buf[29].Feature_n = FeatureBuf_225;
         Mult_Buf[29].Weight_n = Wgt_7_225;
         Mult_Buf[30].Feature_n = FeatureBuf_226;
         Mult_Buf[30].Weight_n = Wgt_7_226;
         Mult_Buf[31].Feature_n = FeatureBuf_227;
         Mult_Buf[31].Weight_n = Wgt_7_227;
         Mult_Buf[32].Feature_n = FeatureBuf_228;
         Mult_Buf[32].Weight_n = Wgt_7_228;
         Mult_Buf[33].Feature_n = FeatureBuf_229;
         Mult_Buf[33].Weight_n = Wgt_7_229;
         Mult_Buf[34].Feature_n = FeatureBuf_230;
         Mult_Buf[34].Weight_n = Wgt_7_230;
         Mult_Buf[35].Feature_n = FeatureBuf_231;
         Mult_Buf[35].Weight_n = Wgt_7_231;
         Mult_Buf[36].Feature_n = FeatureBuf_232;
         Mult_Buf[36].Weight_n = Wgt_7_232;
         Mult_Buf[37].Feature_n = FeatureBuf_233;
         Mult_Buf[37].Weight_n = Wgt_7_233;
         Mult_Buf[38].Feature_n = FeatureBuf_234;
         Mult_Buf[38].Weight_n = Wgt_7_234;
         Mult_Buf[39].Feature_n = FeatureBuf_235;
         Mult_Buf[39].Weight_n = Wgt_7_235;
         Mult_Buf[40].Feature_n = FeatureBuf_236;
         Mult_Buf[40].Weight_n = Wgt_7_236;
         Mult_Buf[41].Feature_n = FeatureBuf_237;
         Mult_Buf[41].Weight_n = Wgt_7_237;
         Mult_Buf[42].Feature_n = FeatureBuf_238;
         Mult_Buf[42].Weight_n = Wgt_7_238;
         Mult_Buf[43].Feature_n = FeatureBuf_239;
         Mult_Buf[43].Weight_n = Wgt_7_239;
         Mult_Buf[44].Feature_n = FeatureBuf_240;
         Mult_Buf[44].Weight_n = Wgt_7_240;
         Mult_Buf[45].Feature_n = FeatureBuf_241;
         Mult_Buf[45].Weight_n = Wgt_7_241;
         Mult_Buf[46].Feature_n = FeatureBuf_242;
         Mult_Buf[46].Weight_n = Wgt_7_242;
         Mult_Buf[47].Feature_n = FeatureBuf_243;
         Mult_Buf[47].Weight_n = Wgt_7_243;
         Mult_Buf[48].Feature_n = FeatureBuf_244;
         Mult_Buf[48].Weight_n = Wgt_7_244;
         Mult_Buf[49].Feature_n = FeatureBuf_245;
         Mult_Buf[49].Weight_n = Wgt_7_245;
         Mult_Buf[50].Feature_n = FeatureBuf_246;
         Mult_Buf[50].Weight_n = Wgt_7_246;
         Mult_Buf[51].Feature_n = FeatureBuf_247;
         Mult_Buf[51].Weight_n = Wgt_7_247;
         Mult_Buf[52].Feature_n = FeatureBuf_248;
         Mult_Buf[52].Weight_n = Wgt_7_248;
         Mult_Buf[53].Feature_n = FeatureBuf_249;
         Mult_Buf[53].Weight_n = Wgt_7_249;
         Mult_Buf[54].Feature_n = FeatureBuf_250;
         Mult_Buf[54].Weight_n = Wgt_7_250;
         Mult_Buf[55].Feature_n = FeatureBuf_251;
         Mult_Buf[55].Weight_n = Wgt_7_251;
         Mult_Buf[56].Feature_n = FeatureBuf_252;
         Mult_Buf[56].Weight_n = Wgt_7_252;
         Mult_Buf[57].Feature_n = FeatureBuf_253;
         Mult_Buf[57].Weight_n = Wgt_7_253;
         Mult_Buf[58].Feature_n = FeatureBuf_254;
         Mult_Buf[58].Weight_n = Wgt_7_254;
         Mult_Buf[59].Feature_n = FeatureBuf_255;
         Mult_Buf[59].Weight_n = Wgt_7_255;
         Mult_Buf[60].Feature_n = FeatureBuf_256;
         Mult_Buf[60].Weight_n = Wgt_7_256;
         Mult_Buf[61].Feature_n = FeatureBuf_257;
         Mult_Buf[61].Weight_n = Wgt_7_257;
         Mult_Buf[62].Feature_n = FeatureBuf_258;
         Mult_Buf[62].Weight_n = Wgt_7_258;
         Mult_Buf[63].Feature_n = FeatureBuf_259;
         Mult_Buf[63].Weight_n = Wgt_7_259;
         Mult_Buf[64].Feature_n = FeatureBuf_260;
         Mult_Buf[64].Weight_n = Wgt_7_260;
         Mult_Buf[65].Feature_n = FeatureBuf_261;
         Mult_Buf[65].Weight_n = Wgt_7_261;
         Mult_Buf[66].Feature_n = FeatureBuf_262;
         Mult_Buf[66].Weight_n = Wgt_7_262;
         Mult_Buf[67].Feature_n = FeatureBuf_263;
         Mult_Buf[67].Weight_n = Wgt_7_263;
         Mult_Buf[68].Feature_n = FeatureBuf_264;
         Mult_Buf[68].Weight_n = Wgt_7_264;
         Mult_Buf[69].Feature_n = FeatureBuf_265;
         Mult_Buf[69].Weight_n = Wgt_7_265;
         Mult_Buf[70].Feature_n = FeatureBuf_266;
         Mult_Buf[70].Weight_n = Wgt_7_266;
         Mult_Buf[71].Feature_n = FeatureBuf_267;
         Mult_Buf[71].Weight_n = Wgt_7_267;
         Mult_Buf[72].Feature_n = FeatureBuf_268;
         Mult_Buf[72].Weight_n = Wgt_7_268;
         Mult_Buf[73].Feature_n = FeatureBuf_269;
         Mult_Buf[73].Weight_n = Wgt_7_269;
         Mult_Buf[74].Feature_n = FeatureBuf_270;
         Mult_Buf[74].Weight_n = Wgt_7_270;
         Mult_Buf[75].Feature_n = FeatureBuf_271;
         Mult_Buf[75].Weight_n = Wgt_7_271;
         Mult_Buf[76].Feature_n = FeatureBuf_272;
         Mult_Buf[76].Weight_n = Wgt_7_272;
         Mult_Buf[77].Feature_n = FeatureBuf_273;
         Mult_Buf[77].Weight_n = Wgt_7_273;
         Mult_Buf[78].Feature_n = FeatureBuf_274;
         Mult_Buf[78].Weight_n = Wgt_7_274;
         Mult_Buf[79].Feature_n = FeatureBuf_275;
         Mult_Buf[79].Weight_n = Wgt_7_275;
         Mult_Buf[80].Feature_n = FeatureBuf_276;
         Mult_Buf[80].Weight_n = Wgt_7_276;
         Mult_Buf[81].Feature_n = FeatureBuf_277;
         Mult_Buf[81].Weight_n = Wgt_7_277;
         Mult_Buf[82].Feature_n = FeatureBuf_278;
         Mult_Buf[82].Weight_n = Wgt_7_278;
         Mult_Buf[83].Feature_n = FeatureBuf_279;
         Mult_Buf[83].Weight_n = Wgt_7_279;
         Mult_Buf[84].Feature_n = FeatureBuf_280;
         Mult_Buf[84].Weight_n = Wgt_7_280;
         Mult_Buf[85].Feature_n = FeatureBuf_281;
         Mult_Buf[85].Weight_n = Wgt_7_281;
         Mult_Buf[86].Feature_n = FeatureBuf_282;
         Mult_Buf[86].Weight_n = Wgt_7_282;
         Mult_Buf[87].Feature_n = FeatureBuf_283;
         Mult_Buf[87].Weight_n = Wgt_7_283;
         Mult_Buf[88].Feature_n = FeatureBuf_284;
         Mult_Buf[88].Weight_n = Wgt_7_284;
         Mult_Buf[89].Feature_n = FeatureBuf_285;
         Mult_Buf[89].Weight_n = Wgt_7_285;
         Mult_Buf[90].Feature_n = FeatureBuf_286;
         Mult_Buf[90].Weight_n = Wgt_7_286;
         Mult_Buf[91].Feature_n = FeatureBuf_287;
         Mult_Buf[91].Weight_n = Wgt_7_287;
         Mult_Buf[92].Feature_n = FeatureBuf_288;
         Mult_Buf[92].Weight_n = Wgt_7_288;
         Mult_Buf[93].Feature_n = FeatureBuf_289;
         Mult_Buf[93].Weight_n = Wgt_7_289;
         Mult_Buf[94].Feature_n = FeatureBuf_290;
         Mult_Buf[94].Weight_n = Wgt_7_290;
         Mult_Buf[95].Feature_n = FeatureBuf_291;
         Mult_Buf[95].Weight_n = Wgt_7_291;
         Mult_Buf[96].Feature_n = FeatureBuf_292;
         Mult_Buf[96].Weight_n = Wgt_7_292;
         Mult_Buf[97].Feature_n = FeatureBuf_293;
         Mult_Buf[97].Weight_n = Wgt_7_293;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     //Collect Partial result form Adder
         Res_4_4_n = Part_Res;
     end
    61:begin
     nxt_state = 62;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_294;
         Mult_Buf[0].Weight_n = Wgt_7_294;
         Mult_Buf[1].Feature_n = FeatureBuf_295;
         Mult_Buf[1].Weight_n = Wgt_7_295;
         Mult_Buf[2].Feature_n = FeatureBuf_296;
         Mult_Buf[2].Weight_n = Wgt_7_296;
         Mult_Buf[3].Feature_n = FeatureBuf_297;
         Mult_Buf[3].Weight_n = Wgt_7_297;
         Mult_Buf[4].Feature_n = FeatureBuf_298;
         Mult_Buf[4].Weight_n = Wgt_7_298;
         Mult_Buf[5].Feature_n = FeatureBuf_299;
         Mult_Buf[5].Weight_n = Wgt_7_299;
         Mult_Buf[6].Feature_n = FeatureBuf_300;
         Mult_Buf[6].Weight_n = Wgt_7_300;
         Mult_Buf[7].Feature_n = FeatureBuf_301;
         Mult_Buf[7].Weight_n = Wgt_7_301;
         Mult_Buf[8].Feature_n = FeatureBuf_302;
         Mult_Buf[8].Weight_n = Wgt_7_302;
         Mult_Buf[9].Feature_n = FeatureBuf_303;
         Mult_Buf[9].Weight_n = Wgt_7_303;
         Mult_Buf[10].Feature_n = FeatureBuf_304;
         Mult_Buf[10].Weight_n = Wgt_7_304;
         Mult_Buf[11].Feature_n = FeatureBuf_305;
         Mult_Buf[11].Weight_n = Wgt_7_305;
         Mult_Buf[12].Feature_n = FeatureBuf_306;
         Mult_Buf[12].Weight_n = Wgt_7_306;
         Mult_Buf[13].Feature_n = FeatureBuf_307;
         Mult_Buf[13].Weight_n = Wgt_7_307;
         Mult_Buf[14].Feature_n = FeatureBuf_308;
         Mult_Buf[14].Weight_n = Wgt_7_308;
         Mult_Buf[15].Feature_n = FeatureBuf_309;
         Mult_Buf[15].Weight_n = Wgt_7_309;
         Mult_Buf[16].Feature_n = FeatureBuf_310;
         Mult_Buf[16].Weight_n = Wgt_7_310;
         Mult_Buf[17].Feature_n = FeatureBuf_311;
         Mult_Buf[17].Weight_n = Wgt_7_311;
         Mult_Buf[18].Feature_n = FeatureBuf_312;
         Mult_Buf[18].Weight_n = Wgt_7_312;
         Mult_Buf[19].Feature_n = FeatureBuf_313;
         Mult_Buf[19].Weight_n = Wgt_7_313;
         Mult_Buf[20].Feature_n = FeatureBuf_314;
         Mult_Buf[20].Weight_n = Wgt_7_314;
         Mult_Buf[21].Feature_n = FeatureBuf_315;
         Mult_Buf[21].Weight_n = Wgt_7_315;
         Mult_Buf[22].Feature_n = FeatureBuf_316;
         Mult_Buf[22].Weight_n = Wgt_7_316;
         Mult_Buf[23].Feature_n = FeatureBuf_317;
         Mult_Buf[23].Weight_n = Wgt_7_317;
         Mult_Buf[24].Feature_n = FeatureBuf_318;
         Mult_Buf[24].Weight_n = Wgt_7_318;
         Mult_Buf[25].Feature_n = FeatureBuf_319;
         Mult_Buf[25].Weight_n = Wgt_7_319;
         Mult_Buf[26].Feature_n = FeatureBuf_320;
         Mult_Buf[26].Weight_n = Wgt_7_320;
         Mult_Buf[27].Feature_n = FeatureBuf_321;
         Mult_Buf[27].Weight_n = Wgt_7_321;
         Mult_Buf[28].Feature_n = FeatureBuf_322;
         Mult_Buf[28].Weight_n = Wgt_7_322;
         Mult_Buf[29].Feature_n = FeatureBuf_323;
         Mult_Buf[29].Weight_n = Wgt_7_323;
         Mult_Buf[30].Feature_n = FeatureBuf_324;
         Mult_Buf[30].Weight_n = Wgt_7_324;
         Mult_Buf[31].Feature_n = FeatureBuf_325;
         Mult_Buf[31].Weight_n = Wgt_7_325;
         Mult_Buf[32].Feature_n = FeatureBuf_326;
         Mult_Buf[32].Weight_n = Wgt_7_326;
         Mult_Buf[33].Feature_n = FeatureBuf_327;
         Mult_Buf[33].Weight_n = Wgt_7_327;
         Mult_Buf[34].Feature_n = FeatureBuf_328;
         Mult_Buf[34].Weight_n = Wgt_7_328;
         Mult_Buf[35].Feature_n = FeatureBuf_329;
         Mult_Buf[35].Weight_n = Wgt_7_329;
         Mult_Buf[36].Feature_n = FeatureBuf_330;
         Mult_Buf[36].Weight_n = Wgt_7_330;
         Mult_Buf[37].Feature_n = FeatureBuf_331;
         Mult_Buf[37].Weight_n = Wgt_7_331;
         Mult_Buf[38].Feature_n = FeatureBuf_332;
         Mult_Buf[38].Weight_n = Wgt_7_332;
         Mult_Buf[39].Feature_n = FeatureBuf_333;
         Mult_Buf[39].Weight_n = Wgt_7_333;
         Mult_Buf[40].Feature_n = FeatureBuf_334;
         Mult_Buf[40].Weight_n = Wgt_7_334;
         Mult_Buf[41].Feature_n = FeatureBuf_335;
         Mult_Buf[41].Weight_n = Wgt_7_335;
         Mult_Buf[42].Feature_n = FeatureBuf_336;
         Mult_Buf[42].Weight_n = Wgt_7_336;
         Mult_Buf[43].Feature_n = FeatureBuf_337;
         Mult_Buf[43].Weight_n = Wgt_7_337;
         Mult_Buf[44].Feature_n = FeatureBuf_338;
         Mult_Buf[44].Weight_n = Wgt_7_338;
         Mult_Buf[45].Feature_n = FeatureBuf_339;
         Mult_Buf[45].Weight_n = Wgt_7_339;
         Mult_Buf[46].Feature_n = FeatureBuf_340;
         Mult_Buf[46].Weight_n = Wgt_7_340;
         Mult_Buf[47].Feature_n = FeatureBuf_341;
         Mult_Buf[47].Weight_n = Wgt_7_341;
         Mult_Buf[48].Feature_n = FeatureBuf_342;
         Mult_Buf[48].Weight_n = Wgt_7_342;
         Mult_Buf[49].Feature_n = FeatureBuf_343;
         Mult_Buf[49].Weight_n = Wgt_7_343;
         Mult_Buf[50].Feature_n = FeatureBuf_344;
         Mult_Buf[50].Weight_n = Wgt_7_344;
         Mult_Buf[51].Feature_n = FeatureBuf_345;
         Mult_Buf[51].Weight_n = Wgt_7_345;
         Mult_Buf[52].Feature_n = FeatureBuf_346;
         Mult_Buf[52].Weight_n = Wgt_7_346;
         Mult_Buf[53].Feature_n = FeatureBuf_347;
         Mult_Buf[53].Weight_n = Wgt_7_347;
         Mult_Buf[54].Feature_n = FeatureBuf_348;
         Mult_Buf[54].Weight_n = Wgt_7_348;
         Mult_Buf[55].Feature_n = FeatureBuf_349;
         Mult_Buf[55].Weight_n = Wgt_7_349;
         Mult_Buf[56].Feature_n = FeatureBuf_350;
         Mult_Buf[56].Weight_n = Wgt_7_350;
         Mult_Buf[57].Feature_n = FeatureBuf_351;
         Mult_Buf[57].Weight_n = Wgt_7_351;
         Mult_Buf[58].Feature_n = FeatureBuf_352;
         Mult_Buf[58].Weight_n = Wgt_7_352;
         Mult_Buf[59].Feature_n = FeatureBuf_353;
         Mult_Buf[59].Weight_n = Wgt_7_353;
         Mult_Buf[60].Feature_n = FeatureBuf_354;
         Mult_Buf[60].Weight_n = Wgt_7_354;
         Mult_Buf[61].Feature_n = FeatureBuf_355;
         Mult_Buf[61].Weight_n = Wgt_7_355;
         Mult_Buf[62].Feature_n = FeatureBuf_356;
         Mult_Buf[62].Weight_n = Wgt_7_356;
         Mult_Buf[63].Feature_n = FeatureBuf_357;
         Mult_Buf[63].Weight_n = Wgt_7_357;
         Mult_Buf[64].Feature_n = FeatureBuf_358;
         Mult_Buf[64].Weight_n = Wgt_7_358;
         Mult_Buf[65].Feature_n = FeatureBuf_359;
         Mult_Buf[65].Weight_n = Wgt_7_359;
         Mult_Buf[66].Feature_n = FeatureBuf_360;
         Mult_Buf[66].Weight_n = Wgt_7_360;
         Mult_Buf[67].Feature_n = FeatureBuf_361;
         Mult_Buf[67].Weight_n = Wgt_7_361;
         Mult_Buf[68].Feature_n = FeatureBuf_362;
         Mult_Buf[68].Weight_n = Wgt_7_362;
         Mult_Buf[69].Feature_n = FeatureBuf_363;
         Mult_Buf[69].Weight_n = Wgt_7_363;
         Mult_Buf[70].Feature_n = FeatureBuf_364;
         Mult_Buf[70].Weight_n = Wgt_7_364;
         Mult_Buf[71].Feature_n = FeatureBuf_365;
         Mult_Buf[71].Weight_n = Wgt_7_365;
         Mult_Buf[72].Feature_n = FeatureBuf_366;
         Mult_Buf[72].Weight_n = Wgt_7_366;
         Mult_Buf[73].Feature_n = FeatureBuf_367;
         Mult_Buf[73].Weight_n = Wgt_7_367;
         Mult_Buf[74].Feature_n = FeatureBuf_368;
         Mult_Buf[74].Weight_n = Wgt_7_368;
         Mult_Buf[75].Feature_n = FeatureBuf_369;
         Mult_Buf[75].Weight_n = Wgt_7_369;
         Mult_Buf[76].Feature_n = FeatureBuf_370;
         Mult_Buf[76].Weight_n = Wgt_7_370;
         Mult_Buf[77].Feature_n = FeatureBuf_371;
         Mult_Buf[77].Weight_n = Wgt_7_371;
         Mult_Buf[78].Feature_n = FeatureBuf_372;
         Mult_Buf[78].Weight_n = Wgt_7_372;
         Mult_Buf[79].Feature_n = FeatureBuf_373;
         Mult_Buf[79].Weight_n = Wgt_7_373;
         Mult_Buf[80].Feature_n = FeatureBuf_374;
         Mult_Buf[80].Weight_n = Wgt_7_374;
         Mult_Buf[81].Feature_n = FeatureBuf_375;
         Mult_Buf[81].Weight_n = Wgt_7_375;
         Mult_Buf[82].Feature_n = FeatureBuf_376;
         Mult_Buf[82].Weight_n = Wgt_7_376;
         Mult_Buf[83].Feature_n = FeatureBuf_377;
         Mult_Buf[83].Weight_n = Wgt_7_377;
         Mult_Buf[84].Feature_n = FeatureBuf_378;
         Mult_Buf[84].Weight_n = Wgt_7_378;
         Mult_Buf[85].Feature_n = FeatureBuf_379;
         Mult_Buf[85].Weight_n = Wgt_7_379;
         Mult_Buf[86].Feature_n = FeatureBuf_380;
         Mult_Buf[86].Weight_n = Wgt_7_380;
         Mult_Buf[87].Feature_n = FeatureBuf_381;
         Mult_Buf[87].Weight_n = Wgt_7_381;
         Mult_Buf[88].Feature_n = FeatureBuf_382;
         Mult_Buf[88].Weight_n = Wgt_7_382;
         Mult_Buf[89].Feature_n = FeatureBuf_383;
         Mult_Buf[89].Weight_n = Wgt_7_383;
         Mult_Buf[90].Feature_n = FeatureBuf_384;
         Mult_Buf[90].Weight_n = Wgt_7_384;
         Mult_Buf[91].Feature_n = FeatureBuf_385;
         Mult_Buf[91].Weight_n = Wgt_7_385;
         Mult_Buf[92].Feature_n = FeatureBuf_386;
         Mult_Buf[92].Weight_n = Wgt_7_386;
         Mult_Buf[93].Feature_n = FeatureBuf_387;
         Mult_Buf[93].Weight_n = Wgt_7_387;
         Mult_Buf[94].Feature_n = FeatureBuf_388;
         Mult_Buf[94].Weight_n = Wgt_7_388;
         Mult_Buf[95].Feature_n = FeatureBuf_389;
         Mult_Buf[95].Weight_n = Wgt_7_389;
         Mult_Buf[96].Feature_n = FeatureBuf_390;
         Mult_Buf[96].Weight_n = Wgt_7_390;
         Mult_Buf[97].Feature_n = FeatureBuf_391;
         Mult_Buf[97].Weight_n = Wgt_7_391;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     //Collect Partial result form Adder
         Res_4_5_n = Part_Res;
     //Collect result from final Adder
         Res3_n = Final_Res;
     end
    62:begin
     nxt_state = 63;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_392;
         Mult_Buf[0].Weight_n = Wgt_7_392;
         Mult_Buf[1].Feature_n = FeatureBuf_393;
         Mult_Buf[1].Weight_n = Wgt_7_393;
         Mult_Buf[2].Feature_n = FeatureBuf_394;
         Mult_Buf[2].Weight_n = Wgt_7_394;
         Mult_Buf[3].Feature_n = FeatureBuf_395;
         Mult_Buf[3].Weight_n = Wgt_7_395;
         Mult_Buf[4].Feature_n = FeatureBuf_396;
         Mult_Buf[4].Weight_n = Wgt_7_396;
         Mult_Buf[5].Feature_n = FeatureBuf_397;
         Mult_Buf[5].Weight_n = Wgt_7_397;
         Mult_Buf[6].Feature_n = FeatureBuf_398;
         Mult_Buf[6].Weight_n = Wgt_7_398;
         Mult_Buf[7].Feature_n = FeatureBuf_399;
         Mult_Buf[7].Weight_n = Wgt_7_399;
         Mult_Buf[8].Feature_n = FeatureBuf_400;
         Mult_Buf[8].Weight_n = Wgt_7_400;
         Mult_Buf[9].Feature_n = FeatureBuf_401;
         Mult_Buf[9].Weight_n = Wgt_7_401;
         Mult_Buf[10].Feature_n = FeatureBuf_402;
         Mult_Buf[10].Weight_n = Wgt_7_402;
         Mult_Buf[11].Feature_n = FeatureBuf_403;
         Mult_Buf[11].Weight_n = Wgt_7_403;
         Mult_Buf[12].Feature_n = FeatureBuf_404;
         Mult_Buf[12].Weight_n = Wgt_7_404;
         Mult_Buf[13].Feature_n = FeatureBuf_405;
         Mult_Buf[13].Weight_n = Wgt_7_405;
         Mult_Buf[14].Feature_n = FeatureBuf_406;
         Mult_Buf[14].Weight_n = Wgt_7_406;
         Mult_Buf[15].Feature_n = FeatureBuf_407;
         Mult_Buf[15].Weight_n = Wgt_7_407;
         Mult_Buf[16].Feature_n = FeatureBuf_408;
         Mult_Buf[16].Weight_n = Wgt_7_408;
         Mult_Buf[17].Feature_n = FeatureBuf_409;
         Mult_Buf[17].Weight_n = Wgt_7_409;
         Mult_Buf[18].Feature_n = FeatureBuf_410;
         Mult_Buf[18].Weight_n = Wgt_7_410;
         Mult_Buf[19].Feature_n = FeatureBuf_411;
         Mult_Buf[19].Weight_n = Wgt_7_411;
         Mult_Buf[20].Feature_n = FeatureBuf_412;
         Mult_Buf[20].Weight_n = Wgt_7_412;
         Mult_Buf[21].Feature_n = FeatureBuf_413;
         Mult_Buf[21].Weight_n = Wgt_7_413;
         Mult_Buf[22].Feature_n = FeatureBuf_414;
         Mult_Buf[22].Weight_n = Wgt_7_414;
         Mult_Buf[23].Feature_n = FeatureBuf_415;
         Mult_Buf[23].Weight_n = Wgt_7_415;
         Mult_Buf[24].Feature_n = FeatureBuf_416;
         Mult_Buf[24].Weight_n = Wgt_7_416;
         Mult_Buf[25].Feature_n = FeatureBuf_417;
         Mult_Buf[25].Weight_n = Wgt_7_417;
         Mult_Buf[26].Feature_n = FeatureBuf_418;
         Mult_Buf[26].Weight_n = Wgt_7_418;
         Mult_Buf[27].Feature_n = FeatureBuf_419;
         Mult_Buf[27].Weight_n = Wgt_7_419;
         Mult_Buf[28].Feature_n = FeatureBuf_420;
         Mult_Buf[28].Weight_n = Wgt_7_420;
         Mult_Buf[29].Feature_n = FeatureBuf_421;
         Mult_Buf[29].Weight_n = Wgt_7_421;
         Mult_Buf[30].Feature_n = FeatureBuf_422;
         Mult_Buf[30].Weight_n = Wgt_7_422;
         Mult_Buf[31].Feature_n = FeatureBuf_423;
         Mult_Buf[31].Weight_n = Wgt_7_423;
         Mult_Buf[32].Feature_n = FeatureBuf_424;
         Mult_Buf[32].Weight_n = Wgt_7_424;
         Mult_Buf[33].Feature_n = FeatureBuf_425;
         Mult_Buf[33].Weight_n = Wgt_7_425;
         Mult_Buf[34].Feature_n = FeatureBuf_426;
         Mult_Buf[34].Weight_n = Wgt_7_426;
         Mult_Buf[35].Feature_n = FeatureBuf_427;
         Mult_Buf[35].Weight_n = Wgt_7_427;
         Mult_Buf[36].Feature_n = FeatureBuf_428;
         Mult_Buf[36].Weight_n = Wgt_7_428;
         Mult_Buf[37].Feature_n = FeatureBuf_429;
         Mult_Buf[37].Weight_n = Wgt_7_429;
         Mult_Buf[38].Feature_n = FeatureBuf_430;
         Mult_Buf[38].Weight_n = Wgt_7_430;
         Mult_Buf[39].Feature_n = FeatureBuf_431;
         Mult_Buf[39].Weight_n = Wgt_7_431;
         Mult_Buf[40].Feature_n = FeatureBuf_432;
         Mult_Buf[40].Weight_n = Wgt_7_432;
         Mult_Buf[41].Feature_n = FeatureBuf_433;
         Mult_Buf[41].Weight_n = Wgt_7_433;
         Mult_Buf[42].Feature_n = FeatureBuf_434;
         Mult_Buf[42].Weight_n = Wgt_7_434;
         Mult_Buf[43].Feature_n = FeatureBuf_435;
         Mult_Buf[43].Weight_n = Wgt_7_435;
         Mult_Buf[44].Feature_n = FeatureBuf_436;
         Mult_Buf[44].Weight_n = Wgt_7_436;
         Mult_Buf[45].Feature_n = FeatureBuf_437;
         Mult_Buf[45].Weight_n = Wgt_7_437;
         Mult_Buf[46].Feature_n = FeatureBuf_438;
         Mult_Buf[46].Weight_n = Wgt_7_438;
         Mult_Buf[47].Feature_n = FeatureBuf_439;
         Mult_Buf[47].Weight_n = Wgt_7_439;
         Mult_Buf[48].Feature_n = FeatureBuf_440;
         Mult_Buf[48].Weight_n = Wgt_7_440;
         Mult_Buf[49].Feature_n = FeatureBuf_441;
         Mult_Buf[49].Weight_n = Wgt_7_441;
         Mult_Buf[50].Feature_n = FeatureBuf_442;
         Mult_Buf[50].Weight_n = Wgt_7_442;
         Mult_Buf[51].Feature_n = FeatureBuf_443;
         Mult_Buf[51].Weight_n = Wgt_7_443;
         Mult_Buf[52].Feature_n = FeatureBuf_444;
         Mult_Buf[52].Weight_n = Wgt_7_444;
         Mult_Buf[53].Feature_n = FeatureBuf_445;
         Mult_Buf[53].Weight_n = Wgt_7_445;
         Mult_Buf[54].Feature_n = FeatureBuf_446;
         Mult_Buf[54].Weight_n = Wgt_7_446;
         Mult_Buf[55].Feature_n = FeatureBuf_447;
         Mult_Buf[55].Weight_n = Wgt_7_447;
         Mult_Buf[56].Feature_n = FeatureBuf_448;
         Mult_Buf[56].Weight_n = Wgt_7_448;
         Mult_Buf[57].Feature_n = FeatureBuf_449;
         Mult_Buf[57].Weight_n = Wgt_7_449;
         Mult_Buf[58].Feature_n = FeatureBuf_450;
         Mult_Buf[58].Weight_n = Wgt_7_450;
         Mult_Buf[59].Feature_n = FeatureBuf_451;
         Mult_Buf[59].Weight_n = Wgt_7_451;
         Mult_Buf[60].Feature_n = FeatureBuf_452;
         Mult_Buf[60].Weight_n = Wgt_7_452;
         Mult_Buf[61].Feature_n = FeatureBuf_453;
         Mult_Buf[61].Weight_n = Wgt_7_453;
         Mult_Buf[62].Feature_n = FeatureBuf_454;
         Mult_Buf[62].Weight_n = Wgt_7_454;
         Mult_Buf[63].Feature_n = FeatureBuf_455;
         Mult_Buf[63].Weight_n = Wgt_7_455;
         Mult_Buf[64].Feature_n = FeatureBuf_456;
         Mult_Buf[64].Weight_n = Wgt_7_456;
         Mult_Buf[65].Feature_n = FeatureBuf_457;
         Mult_Buf[65].Weight_n = Wgt_7_457;
         Mult_Buf[66].Feature_n = FeatureBuf_458;
         Mult_Buf[66].Weight_n = Wgt_7_458;
         Mult_Buf[67].Feature_n = FeatureBuf_459;
         Mult_Buf[67].Weight_n = Wgt_7_459;
         Mult_Buf[68].Feature_n = FeatureBuf_460;
         Mult_Buf[68].Weight_n = Wgt_7_460;
         Mult_Buf[69].Feature_n = FeatureBuf_461;
         Mult_Buf[69].Weight_n = Wgt_7_461;
         Mult_Buf[70].Feature_n = FeatureBuf_462;
         Mult_Buf[70].Weight_n = Wgt_7_462;
         Mult_Buf[71].Feature_n = FeatureBuf_463;
         Mult_Buf[71].Weight_n = Wgt_7_463;
         Mult_Buf[72].Feature_n = FeatureBuf_464;
         Mult_Buf[72].Weight_n = Wgt_7_464;
         Mult_Buf[73].Feature_n = FeatureBuf_465;
         Mult_Buf[73].Weight_n = Wgt_7_465;
         Mult_Buf[74].Feature_n = FeatureBuf_466;
         Mult_Buf[74].Weight_n = Wgt_7_466;
         Mult_Buf[75].Feature_n = FeatureBuf_467;
         Mult_Buf[75].Weight_n = Wgt_7_467;
         Mult_Buf[76].Feature_n = FeatureBuf_468;
         Mult_Buf[76].Weight_n = Wgt_7_468;
         Mult_Buf[77].Feature_n = FeatureBuf_469;
         Mult_Buf[77].Weight_n = Wgt_7_469;
         Mult_Buf[78].Feature_n = FeatureBuf_470;
         Mult_Buf[78].Weight_n = Wgt_7_470;
         Mult_Buf[79].Feature_n = FeatureBuf_471;
         Mult_Buf[79].Weight_n = Wgt_7_471;
         Mult_Buf[80].Feature_n = FeatureBuf_472;
         Mult_Buf[80].Weight_n = Wgt_7_472;
         Mult_Buf[81].Feature_n = FeatureBuf_473;
         Mult_Buf[81].Weight_n = Wgt_7_473;
         Mult_Buf[82].Feature_n = FeatureBuf_474;
         Mult_Buf[82].Weight_n = Wgt_7_474;
         Mult_Buf[83].Feature_n = FeatureBuf_475;
         Mult_Buf[83].Weight_n = Wgt_7_475;
         Mult_Buf[84].Feature_n = FeatureBuf_476;
         Mult_Buf[84].Weight_n = Wgt_7_476;
         Mult_Buf[85].Feature_n = FeatureBuf_477;
         Mult_Buf[85].Weight_n = Wgt_7_477;
         Mult_Buf[86].Feature_n = FeatureBuf_478;
         Mult_Buf[86].Weight_n = Wgt_7_478;
         Mult_Buf[87].Feature_n = FeatureBuf_479;
         Mult_Buf[87].Weight_n = Wgt_7_479;
         Mult_Buf[88].Feature_n = FeatureBuf_480;
         Mult_Buf[88].Weight_n = Wgt_7_480;
         Mult_Buf[89].Feature_n = FeatureBuf_481;
         Mult_Buf[89].Weight_n = Wgt_7_481;
         Mult_Buf[90].Feature_n = FeatureBuf_482;
         Mult_Buf[90].Weight_n = Wgt_7_482;
         Mult_Buf[91].Feature_n = FeatureBuf_483;
         Mult_Buf[91].Weight_n = Wgt_7_483;
         Mult_Buf[92].Feature_n = FeatureBuf_484;
         Mult_Buf[92].Weight_n = Wgt_7_484;
         Mult_Buf[93].Feature_n = FeatureBuf_485;
         Mult_Buf[93].Weight_n = Wgt_7_485;
         Mult_Buf[94].Feature_n = FeatureBuf_486;
         Mult_Buf[94].Weight_n = Wgt_7_486;
         Mult_Buf[95].Feature_n = FeatureBuf_487;
         Mult_Buf[95].Weight_n = Wgt_7_487;
         Mult_Buf[96].Feature_n = FeatureBuf_488;
         Mult_Buf[96].Weight_n = Wgt_7_488;
         Mult_Buf[97].Feature_n = FeatureBuf_489;
         Mult_Buf[97].Weight_n = Wgt_7_489;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     //Collect Partial result form Adder
         Res_4_6_n = Part_Res;
     end
    63:begin
     nxt_state = 64;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_490;
         Mult_Buf[0].Weight_n = Wgt_7_490;
         Mult_Buf[1].Feature_n = FeatureBuf_491;
         Mult_Buf[1].Weight_n = Wgt_7_491;
         Mult_Buf[2].Feature_n = FeatureBuf_492;
         Mult_Buf[2].Weight_n = Wgt_7_492;
         Mult_Buf[3].Feature_n = FeatureBuf_493;
         Mult_Buf[3].Weight_n = Wgt_7_493;
         Mult_Buf[4].Feature_n = FeatureBuf_494;
         Mult_Buf[4].Weight_n = Wgt_7_494;
         Mult_Buf[5].Feature_n = FeatureBuf_495;
         Mult_Buf[5].Weight_n = Wgt_7_495;
         Mult_Buf[6].Feature_n = FeatureBuf_496;
         Mult_Buf[6].Weight_n = Wgt_7_496;
         Mult_Buf[7].Feature_n = FeatureBuf_497;
         Mult_Buf[7].Weight_n = Wgt_7_497;
         Mult_Buf[8].Feature_n = FeatureBuf_498;
         Mult_Buf[8].Weight_n = Wgt_7_498;
         Mult_Buf[9].Feature_n = FeatureBuf_499;
         Mult_Buf[9].Weight_n = Wgt_7_499;
         Mult_Buf[10].Feature_n = FeatureBuf_500;
         Mult_Buf[10].Weight_n = Wgt_7_500;
         Mult_Buf[11].Feature_n = FeatureBuf_501;
         Mult_Buf[11].Weight_n = Wgt_7_501;
         Mult_Buf[12].Feature_n = FeatureBuf_502;
         Mult_Buf[12].Weight_n = Wgt_7_502;
         Mult_Buf[13].Feature_n = FeatureBuf_503;
         Mult_Buf[13].Weight_n = Wgt_7_503;
         Mult_Buf[14].Feature_n = FeatureBuf_504;
         Mult_Buf[14].Weight_n = Wgt_7_504;
         Mult_Buf[15].Feature_n = FeatureBuf_505;
         Mult_Buf[15].Weight_n = Wgt_7_505;
         Mult_Buf[16].Feature_n = FeatureBuf_506;
         Mult_Buf[16].Weight_n = Wgt_7_506;
         Mult_Buf[17].Feature_n = FeatureBuf_507;
         Mult_Buf[17].Weight_n = Wgt_7_507;
         Mult_Buf[18].Feature_n = FeatureBuf_508;
         Mult_Buf[18].Weight_n = Wgt_7_508;
         Mult_Buf[19].Feature_n = FeatureBuf_509;
         Mult_Buf[19].Weight_n = Wgt_7_509;
         Mult_Buf[20].Feature_n = FeatureBuf_510;
         Mult_Buf[20].Weight_n = Wgt_7_510;
         Mult_Buf[21].Feature_n = FeatureBuf_511;
         Mult_Buf[21].Weight_n = Wgt_7_511;
         Mult_Buf[22].Feature_n = FeatureBuf_512;
         Mult_Buf[22].Weight_n = Wgt_7_512;
         Mult_Buf[23].Feature_n = FeatureBuf_513;
         Mult_Buf[23].Weight_n = Wgt_7_513;
         Mult_Buf[24].Feature_n = FeatureBuf_514;
         Mult_Buf[24].Weight_n = Wgt_7_514;
         Mult_Buf[25].Feature_n = FeatureBuf_515;
         Mult_Buf[25].Weight_n = Wgt_7_515;
         Mult_Buf[26].Feature_n = FeatureBuf_516;
         Mult_Buf[26].Weight_n = Wgt_7_516;
         Mult_Buf[27].Feature_n = FeatureBuf_517;
         Mult_Buf[27].Weight_n = Wgt_7_517;
         Mult_Buf[28].Feature_n = FeatureBuf_518;
         Mult_Buf[28].Weight_n = Wgt_7_518;
         Mult_Buf[29].Feature_n = FeatureBuf_519;
         Mult_Buf[29].Weight_n = Wgt_7_519;
         Mult_Buf[30].Feature_n = FeatureBuf_520;
         Mult_Buf[30].Weight_n = Wgt_7_520;
         Mult_Buf[31].Feature_n = FeatureBuf_521;
         Mult_Buf[31].Weight_n = Wgt_7_521;
         Mult_Buf[32].Feature_n = FeatureBuf_522;
         Mult_Buf[32].Weight_n = Wgt_7_522;
         Mult_Buf[33].Feature_n = FeatureBuf_523;
         Mult_Buf[33].Weight_n = Wgt_7_523;
         Mult_Buf[34].Feature_n = FeatureBuf_524;
         Mult_Buf[34].Weight_n = Wgt_7_524;
         Mult_Buf[35].Feature_n = FeatureBuf_525;
         Mult_Buf[35].Weight_n = Wgt_7_525;
         Mult_Buf[36].Feature_n = FeatureBuf_526;
         Mult_Buf[36].Weight_n = Wgt_7_526;
         Mult_Buf[37].Feature_n = FeatureBuf_527;
         Mult_Buf[37].Weight_n = Wgt_7_527;
         Mult_Buf[38].Feature_n = FeatureBuf_528;
         Mult_Buf[38].Weight_n = Wgt_7_528;
         Mult_Buf[39].Feature_n = FeatureBuf_529;
         Mult_Buf[39].Weight_n = Wgt_7_529;
         Mult_Buf[40].Feature_n = FeatureBuf_530;
         Mult_Buf[40].Weight_n = Wgt_7_530;
         Mult_Buf[41].Feature_n = FeatureBuf_531;
         Mult_Buf[41].Weight_n = Wgt_7_531;
         Mult_Buf[42].Feature_n = FeatureBuf_532;
         Mult_Buf[42].Weight_n = Wgt_7_532;
         Mult_Buf[43].Feature_n = FeatureBuf_533;
         Mult_Buf[43].Weight_n = Wgt_7_533;
         Mult_Buf[44].Feature_n = FeatureBuf_534;
         Mult_Buf[44].Weight_n = Wgt_7_534;
         Mult_Buf[45].Feature_n = FeatureBuf_535;
         Mult_Buf[45].Weight_n = Wgt_7_535;
         Mult_Buf[46].Feature_n = FeatureBuf_536;
         Mult_Buf[46].Weight_n = Wgt_7_536;
         Mult_Buf[47].Feature_n = FeatureBuf_537;
         Mult_Buf[47].Weight_n = Wgt_7_537;
         Mult_Buf[48].Feature_n = FeatureBuf_538;
         Mult_Buf[48].Weight_n = Wgt_7_538;
         Mult_Buf[49].Feature_n = FeatureBuf_539;
         Mult_Buf[49].Weight_n = Wgt_7_539;
         Mult_Buf[50].Feature_n = FeatureBuf_540;
         Mult_Buf[50].Weight_n = Wgt_7_540;
         Mult_Buf[51].Feature_n = FeatureBuf_541;
         Mult_Buf[51].Weight_n = Wgt_7_541;
         Mult_Buf[52].Feature_n = FeatureBuf_542;
         Mult_Buf[52].Weight_n = Wgt_7_542;
         Mult_Buf[53].Feature_n = FeatureBuf_543;
         Mult_Buf[53].Weight_n = Wgt_7_543;
         Mult_Buf[54].Feature_n = FeatureBuf_544;
         Mult_Buf[54].Weight_n = Wgt_7_544;
         Mult_Buf[55].Feature_n = FeatureBuf_545;
         Mult_Buf[55].Weight_n = Wgt_7_545;
         Mult_Buf[56].Feature_n = FeatureBuf_546;
         Mult_Buf[56].Weight_n = Wgt_7_546;
         Mult_Buf[57].Feature_n = FeatureBuf_547;
         Mult_Buf[57].Weight_n = Wgt_7_547;
         Mult_Buf[58].Feature_n = FeatureBuf_548;
         Mult_Buf[58].Weight_n = Wgt_7_548;
         Mult_Buf[59].Feature_n = FeatureBuf_549;
         Mult_Buf[59].Weight_n = Wgt_7_549;
         Mult_Buf[60].Feature_n = FeatureBuf_550;
         Mult_Buf[60].Weight_n = Wgt_7_550;
         Mult_Buf[61].Feature_n = FeatureBuf_551;
         Mult_Buf[61].Weight_n = Wgt_7_551;
         Mult_Buf[62].Feature_n = FeatureBuf_552;
         Mult_Buf[62].Weight_n = Wgt_7_552;
         Mult_Buf[63].Feature_n = FeatureBuf_553;
         Mult_Buf[63].Weight_n = Wgt_7_553;
         Mult_Buf[64].Feature_n = FeatureBuf_554;
         Mult_Buf[64].Weight_n = Wgt_7_554;
         Mult_Buf[65].Feature_n = FeatureBuf_555;
         Mult_Buf[65].Weight_n = Wgt_7_555;
         Mult_Buf[66].Feature_n = FeatureBuf_556;
         Mult_Buf[66].Weight_n = Wgt_7_556;
         Mult_Buf[67].Feature_n = FeatureBuf_557;
         Mult_Buf[67].Weight_n = Wgt_7_557;
         Mult_Buf[68].Feature_n = FeatureBuf_558;
         Mult_Buf[68].Weight_n = Wgt_7_558;
         Mult_Buf[69].Feature_n = FeatureBuf_559;
         Mult_Buf[69].Weight_n = Wgt_7_559;
         Mult_Buf[70].Feature_n = FeatureBuf_560;
         Mult_Buf[70].Weight_n = Wgt_7_560;
         Mult_Buf[71].Feature_n = FeatureBuf_561;
         Mult_Buf[71].Weight_n = Wgt_7_561;
         Mult_Buf[72].Feature_n = FeatureBuf_562;
         Mult_Buf[72].Weight_n = Wgt_7_562;
         Mult_Buf[73].Feature_n = FeatureBuf_563;
         Mult_Buf[73].Weight_n = Wgt_7_563;
         Mult_Buf[74].Feature_n = FeatureBuf_564;
         Mult_Buf[74].Weight_n = Wgt_7_564;
         Mult_Buf[75].Feature_n = FeatureBuf_565;
         Mult_Buf[75].Weight_n = Wgt_7_565;
         Mult_Buf[76].Feature_n = FeatureBuf_566;
         Mult_Buf[76].Weight_n = Wgt_7_566;
         Mult_Buf[77].Feature_n = FeatureBuf_567;
         Mult_Buf[77].Weight_n = Wgt_7_567;
         Mult_Buf[78].Feature_n = FeatureBuf_568;
         Mult_Buf[78].Weight_n = Wgt_7_568;
         Mult_Buf[79].Feature_n = FeatureBuf_569;
         Mult_Buf[79].Weight_n = Wgt_7_569;
         Mult_Buf[80].Feature_n = FeatureBuf_570;
         Mult_Buf[80].Weight_n = Wgt_7_570;
         Mult_Buf[81].Feature_n = FeatureBuf_571;
         Mult_Buf[81].Weight_n = Wgt_7_571;
         Mult_Buf[82].Feature_n = FeatureBuf_572;
         Mult_Buf[82].Weight_n = Wgt_7_572;
         Mult_Buf[83].Feature_n = FeatureBuf_573;
         Mult_Buf[83].Weight_n = Wgt_7_573;
         Mult_Buf[84].Feature_n = FeatureBuf_574;
         Mult_Buf[84].Weight_n = Wgt_7_574;
         Mult_Buf[85].Feature_n = FeatureBuf_575;
         Mult_Buf[85].Weight_n = Wgt_7_575;
         Mult_Buf[86].Feature_n = FeatureBuf_576;
         Mult_Buf[86].Weight_n = Wgt_7_576;
         Mult_Buf[87].Feature_n = FeatureBuf_577;
         Mult_Buf[87].Weight_n = Wgt_7_577;
         Mult_Buf[88].Feature_n = FeatureBuf_578;
         Mult_Buf[88].Weight_n = Wgt_7_578;
         Mult_Buf[89].Feature_n = FeatureBuf_579;
         Mult_Buf[89].Weight_n = Wgt_7_579;
         Mult_Buf[90].Feature_n = FeatureBuf_580;
         Mult_Buf[90].Weight_n = Wgt_7_580;
         Mult_Buf[91].Feature_n = FeatureBuf_581;
         Mult_Buf[91].Weight_n = Wgt_7_581;
         Mult_Buf[92].Feature_n = FeatureBuf_582;
         Mult_Buf[92].Weight_n = Wgt_7_582;
         Mult_Buf[93].Feature_n = FeatureBuf_583;
         Mult_Buf[93].Weight_n = Wgt_7_583;
         Mult_Buf[94].Feature_n = FeatureBuf_584;
         Mult_Buf[94].Weight_n = Wgt_7_584;
         Mult_Buf[95].Feature_n = FeatureBuf_585;
         Mult_Buf[95].Weight_n = Wgt_7_585;
         Mult_Buf[96].Feature_n = FeatureBuf_586;
         Mult_Buf[96].Weight_n = Wgt_7_586;
         Mult_Buf[97].Feature_n = FeatureBuf_587;
         Mult_Buf[97].Weight_n = Wgt_7_587;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     //Collect Partial result form Adder
         Res_4_7_n = Part_Res;
     //Feed to final Adder
         A1 = Part_Res;
         A2 = Res_4_6_n;
         A3 = Res_4_5_n;
         A4 = Res_4_4_n;
         A5 = Res_4_3_n;
         A6 = Res_4_2_n;
         A7 = Res_4_1_n;
         A8 = Res_4_0_n;
     end
    64:begin
     nxt_state = 65;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_588;
         Mult_Buf[0].Weight_n = Wgt_7_588;
         Mult_Buf[1].Feature_n = FeatureBuf_589;
         Mult_Buf[1].Weight_n = Wgt_7_589;
         Mult_Buf[2].Feature_n = FeatureBuf_590;
         Mult_Buf[2].Weight_n = Wgt_7_590;
         Mult_Buf[3].Feature_n = FeatureBuf_591;
         Mult_Buf[3].Weight_n = Wgt_7_591;
         Mult_Buf[4].Feature_n = FeatureBuf_592;
         Mult_Buf[4].Weight_n = Wgt_7_592;
         Mult_Buf[5].Feature_n = FeatureBuf_593;
         Mult_Buf[5].Weight_n = Wgt_7_593;
         Mult_Buf[6].Feature_n = FeatureBuf_594;
         Mult_Buf[6].Weight_n = Wgt_7_594;
         Mult_Buf[7].Feature_n = FeatureBuf_595;
         Mult_Buf[7].Weight_n = Wgt_7_595;
         Mult_Buf[8].Feature_n = FeatureBuf_596;
         Mult_Buf[8].Weight_n = Wgt_7_596;
         Mult_Buf[9].Feature_n = FeatureBuf_597;
         Mult_Buf[9].Weight_n = Wgt_7_597;
         Mult_Buf[10].Feature_n = FeatureBuf_598;
         Mult_Buf[10].Weight_n = Wgt_7_598;
         Mult_Buf[11].Feature_n = FeatureBuf_599;
         Mult_Buf[11].Weight_n = Wgt_7_599;
         Mult_Buf[12].Feature_n = FeatureBuf_600;
         Mult_Buf[12].Weight_n = Wgt_7_600;
         Mult_Buf[13].Feature_n = FeatureBuf_601;
         Mult_Buf[13].Weight_n = Wgt_7_601;
         Mult_Buf[14].Feature_n = FeatureBuf_602;
         Mult_Buf[14].Weight_n = Wgt_7_602;
         Mult_Buf[15].Feature_n = FeatureBuf_603;
         Mult_Buf[15].Weight_n = Wgt_7_603;
         Mult_Buf[16].Feature_n = FeatureBuf_604;
         Mult_Buf[16].Weight_n = Wgt_7_604;
         Mult_Buf[17].Feature_n = FeatureBuf_605;
         Mult_Buf[17].Weight_n = Wgt_7_605;
         Mult_Buf[18].Feature_n = FeatureBuf_606;
         Mult_Buf[18].Weight_n = Wgt_7_606;
         Mult_Buf[19].Feature_n = FeatureBuf_607;
         Mult_Buf[19].Weight_n = Wgt_7_607;
         Mult_Buf[20].Feature_n = FeatureBuf_608;
         Mult_Buf[20].Weight_n = Wgt_7_608;
         Mult_Buf[21].Feature_n = FeatureBuf_609;
         Mult_Buf[21].Weight_n = Wgt_7_609;
         Mult_Buf[22].Feature_n = FeatureBuf_610;
         Mult_Buf[22].Weight_n = Wgt_7_610;
         Mult_Buf[23].Feature_n = FeatureBuf_611;
         Mult_Buf[23].Weight_n = Wgt_7_611;
         Mult_Buf[24].Feature_n = FeatureBuf_612;
         Mult_Buf[24].Weight_n = Wgt_7_612;
         Mult_Buf[25].Feature_n = FeatureBuf_613;
         Mult_Buf[25].Weight_n = Wgt_7_613;
         Mult_Buf[26].Feature_n = FeatureBuf_614;
         Mult_Buf[26].Weight_n = Wgt_7_614;
         Mult_Buf[27].Feature_n = FeatureBuf_615;
         Mult_Buf[27].Weight_n = Wgt_7_615;
         Mult_Buf[28].Feature_n = FeatureBuf_616;
         Mult_Buf[28].Weight_n = Wgt_7_616;
         Mult_Buf[29].Feature_n = FeatureBuf_617;
         Mult_Buf[29].Weight_n = Wgt_7_617;
         Mult_Buf[30].Feature_n = FeatureBuf_618;
         Mult_Buf[30].Weight_n = Wgt_7_618;
         Mult_Buf[31].Feature_n = FeatureBuf_619;
         Mult_Buf[31].Weight_n = Wgt_7_619;
         Mult_Buf[32].Feature_n = FeatureBuf_620;
         Mult_Buf[32].Weight_n = Wgt_7_620;
         Mult_Buf[33].Feature_n = FeatureBuf_621;
         Mult_Buf[33].Weight_n = Wgt_7_621;
         Mult_Buf[34].Feature_n = FeatureBuf_622;
         Mult_Buf[34].Weight_n = Wgt_7_622;
         Mult_Buf[35].Feature_n = FeatureBuf_623;
         Mult_Buf[35].Weight_n = Wgt_7_623;
         Mult_Buf[36].Feature_n = FeatureBuf_624;
         Mult_Buf[36].Weight_n = Wgt_7_624;
         Mult_Buf[37].Feature_n = FeatureBuf_625;
         Mult_Buf[37].Weight_n = Wgt_7_625;
         Mult_Buf[38].Feature_n = FeatureBuf_626;
         Mult_Buf[38].Weight_n = Wgt_7_626;
         Mult_Buf[39].Feature_n = FeatureBuf_627;
         Mult_Buf[39].Weight_n = Wgt_7_627;
         Mult_Buf[40].Feature_n = FeatureBuf_628;
         Mult_Buf[40].Weight_n = Wgt_7_628;
         Mult_Buf[41].Feature_n = FeatureBuf_629;
         Mult_Buf[41].Weight_n = Wgt_7_629;
         Mult_Buf[42].Feature_n = FeatureBuf_630;
         Mult_Buf[42].Weight_n = Wgt_7_630;
         Mult_Buf[43].Feature_n = FeatureBuf_631;
         Mult_Buf[43].Weight_n = Wgt_7_631;
         Mult_Buf[44].Feature_n = FeatureBuf_632;
         Mult_Buf[44].Weight_n = Wgt_7_632;
         Mult_Buf[45].Feature_n = FeatureBuf_633;
         Mult_Buf[45].Weight_n = Wgt_7_633;
         Mult_Buf[46].Feature_n = FeatureBuf_634;
         Mult_Buf[46].Weight_n = Wgt_7_634;
         Mult_Buf[47].Feature_n = FeatureBuf_635;
         Mult_Buf[47].Weight_n = Wgt_7_635;
         Mult_Buf[48].Feature_n = FeatureBuf_636;
         Mult_Buf[48].Weight_n = Wgt_7_636;
         Mult_Buf[49].Feature_n = FeatureBuf_637;
         Mult_Buf[49].Weight_n = Wgt_7_637;
         Mult_Buf[50].Feature_n = FeatureBuf_638;
         Mult_Buf[50].Weight_n = Wgt_7_638;
         Mult_Buf[51].Feature_n = FeatureBuf_639;
         Mult_Buf[51].Weight_n = Wgt_7_639;
         Mult_Buf[52].Feature_n = FeatureBuf_640;
         Mult_Buf[52].Weight_n = Wgt_7_640;
         Mult_Buf[53].Feature_n = FeatureBuf_641;
         Mult_Buf[53].Weight_n = Wgt_7_641;
         Mult_Buf[54].Feature_n = FeatureBuf_642;
         Mult_Buf[54].Weight_n = Wgt_7_642;
         Mult_Buf[55].Feature_n = FeatureBuf_643;
         Mult_Buf[55].Weight_n = Wgt_7_643;
         Mult_Buf[56].Feature_n = FeatureBuf_644;
         Mult_Buf[56].Weight_n = Wgt_7_644;
         Mult_Buf[57].Feature_n = FeatureBuf_645;
         Mult_Buf[57].Weight_n = Wgt_7_645;
         Mult_Buf[58].Feature_n = FeatureBuf_646;
         Mult_Buf[58].Weight_n = Wgt_7_646;
         Mult_Buf[59].Feature_n = FeatureBuf_647;
         Mult_Buf[59].Weight_n = Wgt_7_647;
         Mult_Buf[60].Feature_n = FeatureBuf_648;
         Mult_Buf[60].Weight_n = Wgt_7_648;
         Mult_Buf[61].Feature_n = FeatureBuf_649;
         Mult_Buf[61].Weight_n = Wgt_7_649;
         Mult_Buf[62].Feature_n = FeatureBuf_650;
         Mult_Buf[62].Weight_n = Wgt_7_650;
         Mult_Buf[63].Feature_n = FeatureBuf_651;
         Mult_Buf[63].Weight_n = Wgt_7_651;
         Mult_Buf[64].Feature_n = FeatureBuf_652;
         Mult_Buf[64].Weight_n = Wgt_7_652;
         Mult_Buf[65].Feature_n = FeatureBuf_653;
         Mult_Buf[65].Weight_n = Wgt_7_653;
         Mult_Buf[66].Feature_n = FeatureBuf_654;
         Mult_Buf[66].Weight_n = Wgt_7_654;
         Mult_Buf[67].Feature_n = FeatureBuf_655;
         Mult_Buf[67].Weight_n = Wgt_7_655;
         Mult_Buf[68].Feature_n = FeatureBuf_656;
         Mult_Buf[68].Weight_n = Wgt_7_656;
         Mult_Buf[69].Feature_n = FeatureBuf_657;
         Mult_Buf[69].Weight_n = Wgt_7_657;
         Mult_Buf[70].Feature_n = FeatureBuf_658;
         Mult_Buf[70].Weight_n = Wgt_7_658;
         Mult_Buf[71].Feature_n = FeatureBuf_659;
         Mult_Buf[71].Weight_n = Wgt_7_659;
         Mult_Buf[72].Feature_n = FeatureBuf_660;
         Mult_Buf[72].Weight_n = Wgt_7_660;
         Mult_Buf[73].Feature_n = FeatureBuf_661;
         Mult_Buf[73].Weight_n = Wgt_7_661;
         Mult_Buf[74].Feature_n = FeatureBuf_662;
         Mult_Buf[74].Weight_n = Wgt_7_662;
         Mult_Buf[75].Feature_n = FeatureBuf_663;
         Mult_Buf[75].Weight_n = Wgt_7_663;
         Mult_Buf[76].Feature_n = FeatureBuf_664;
         Mult_Buf[76].Weight_n = Wgt_7_664;
         Mult_Buf[77].Feature_n = FeatureBuf_665;
         Mult_Buf[77].Weight_n = Wgt_7_665;
         Mult_Buf[78].Feature_n = FeatureBuf_666;
         Mult_Buf[78].Weight_n = Wgt_7_666;
         Mult_Buf[79].Feature_n = FeatureBuf_667;
         Mult_Buf[79].Weight_n = Wgt_7_667;
         Mult_Buf[80].Feature_n = FeatureBuf_668;
         Mult_Buf[80].Weight_n = Wgt_7_668;
         Mult_Buf[81].Feature_n = FeatureBuf_669;
         Mult_Buf[81].Weight_n = Wgt_7_669;
         Mult_Buf[82].Feature_n = FeatureBuf_670;
         Mult_Buf[82].Weight_n = Wgt_7_670;
         Mult_Buf[83].Feature_n = FeatureBuf_671;
         Mult_Buf[83].Weight_n = Wgt_7_671;
         Mult_Buf[84].Feature_n = FeatureBuf_672;
         Mult_Buf[84].Weight_n = Wgt_7_672;
         Mult_Buf[85].Feature_n = FeatureBuf_673;
         Mult_Buf[85].Weight_n = Wgt_7_673;
         Mult_Buf[86].Feature_n = FeatureBuf_674;
         Mult_Buf[86].Weight_n = Wgt_7_674;
         Mult_Buf[87].Feature_n = FeatureBuf_675;
         Mult_Buf[87].Weight_n = Wgt_7_675;
         Mult_Buf[88].Feature_n = FeatureBuf_676;
         Mult_Buf[88].Weight_n = Wgt_7_676;
         Mult_Buf[89].Feature_n = FeatureBuf_677;
         Mult_Buf[89].Weight_n = Wgt_7_677;
         Mult_Buf[90].Feature_n = FeatureBuf_678;
         Mult_Buf[90].Weight_n = Wgt_7_678;
         Mult_Buf[91].Feature_n = FeatureBuf_679;
         Mult_Buf[91].Weight_n = Wgt_7_679;
         Mult_Buf[92].Feature_n = FeatureBuf_680;
         Mult_Buf[92].Weight_n = Wgt_7_680;
         Mult_Buf[93].Feature_n = FeatureBuf_681;
         Mult_Buf[93].Weight_n = Wgt_7_681;
         Mult_Buf[94].Feature_n = FeatureBuf_682;
         Mult_Buf[94].Weight_n = Wgt_7_682;
         Mult_Buf[95].Feature_n = FeatureBuf_683;
         Mult_Buf[95].Weight_n = Wgt_7_683;
         Mult_Buf[96].Feature_n = FeatureBuf_684;
         Mult_Buf[96].Weight_n = Wgt_7_684;
         Mult_Buf[97].Feature_n = FeatureBuf_685;
         Mult_Buf[97].Weight_n = Wgt_7_685;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     //Collect Partial result form Adder
         Res_5_0_n = Part_Res;
     end
    65:begin
     nxt_state = 66;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_686;
         Mult_Buf[0].Weight_n = Wgt_7_686;
         Mult_Buf[1].Feature_n = FeatureBuf_687;
         Mult_Buf[1].Weight_n = Wgt_7_687;
         Mult_Buf[2].Feature_n = FeatureBuf_688;
         Mult_Buf[2].Weight_n = Wgt_7_688;
         Mult_Buf[3].Feature_n = FeatureBuf_689;
         Mult_Buf[3].Weight_n = Wgt_7_689;
         Mult_Buf[4].Feature_n = FeatureBuf_690;
         Mult_Buf[4].Weight_n = Wgt_7_690;
         Mult_Buf[5].Feature_n = FeatureBuf_691;
         Mult_Buf[5].Weight_n = Wgt_7_691;
         Mult_Buf[6].Feature_n = FeatureBuf_692;
         Mult_Buf[6].Weight_n = Wgt_7_692;
         Mult_Buf[7].Feature_n = FeatureBuf_693;
         Mult_Buf[7].Weight_n = Wgt_7_693;
         Mult_Buf[8].Feature_n = FeatureBuf_694;
         Mult_Buf[8].Weight_n = Wgt_7_694;
         Mult_Buf[9].Feature_n = FeatureBuf_695;
         Mult_Buf[9].Weight_n = Wgt_7_695;
         Mult_Buf[10].Feature_n = FeatureBuf_696;
         Mult_Buf[10].Weight_n = Wgt_7_696;
         Mult_Buf[11].Feature_n = FeatureBuf_697;
         Mult_Buf[11].Weight_n = Wgt_7_697;
         Mult_Buf[12].Feature_n = FeatureBuf_698;
         Mult_Buf[12].Weight_n = Wgt_7_698;
         Mult_Buf[13].Feature_n = FeatureBuf_699;
         Mult_Buf[13].Weight_n = Wgt_7_699;
         Mult_Buf[14].Feature_n = FeatureBuf_700;
         Mult_Buf[14].Weight_n = Wgt_7_700;
         Mult_Buf[15].Feature_n = FeatureBuf_701;
         Mult_Buf[15].Weight_n = Wgt_7_701;
         Mult_Buf[16].Feature_n = FeatureBuf_702;
         Mult_Buf[16].Weight_n = Wgt_7_702;
         Mult_Buf[17].Feature_n = FeatureBuf_703;
         Mult_Buf[17].Weight_n = Wgt_7_703;
         Mult_Buf[18].Feature_n = FeatureBuf_704;
         Mult_Buf[18].Weight_n = Wgt_7_704;
         Mult_Buf[19].Feature_n = FeatureBuf_705;
         Mult_Buf[19].Weight_n = Wgt_7_705;
         Mult_Buf[20].Feature_n = FeatureBuf_706;
         Mult_Buf[20].Weight_n = Wgt_7_706;
         Mult_Buf[21].Feature_n = FeatureBuf_707;
         Mult_Buf[21].Weight_n = Wgt_7_707;
         Mult_Buf[22].Feature_n = FeatureBuf_708;
         Mult_Buf[22].Weight_n = Wgt_7_708;
         Mult_Buf[23].Feature_n = FeatureBuf_709;
         Mult_Buf[23].Weight_n = Wgt_7_709;
         Mult_Buf[24].Feature_n = FeatureBuf_710;
         Mult_Buf[24].Weight_n = Wgt_7_710;
         Mult_Buf[25].Feature_n = FeatureBuf_711;
         Mult_Buf[25].Weight_n = Wgt_7_711;
         Mult_Buf[26].Feature_n = FeatureBuf_712;
         Mult_Buf[26].Weight_n = Wgt_7_712;
         Mult_Buf[27].Feature_n = FeatureBuf_713;
         Mult_Buf[27].Weight_n = Wgt_7_713;
         Mult_Buf[28].Feature_n = FeatureBuf_714;
         Mult_Buf[28].Weight_n = Wgt_7_714;
         Mult_Buf[29].Feature_n = FeatureBuf_715;
         Mult_Buf[29].Weight_n = Wgt_7_715;
         Mult_Buf[30].Feature_n = FeatureBuf_716;
         Mult_Buf[30].Weight_n = Wgt_7_716;
         Mult_Buf[31].Feature_n = FeatureBuf_717;
         Mult_Buf[31].Weight_n = Wgt_7_717;
         Mult_Buf[32].Feature_n = FeatureBuf_718;
         Mult_Buf[32].Weight_n = Wgt_7_718;
         Mult_Buf[33].Feature_n = FeatureBuf_719;
         Mult_Buf[33].Weight_n = Wgt_7_719;
         Mult_Buf[34].Feature_n = FeatureBuf_720;
         Mult_Buf[34].Weight_n = Wgt_7_720;
         Mult_Buf[35].Feature_n = FeatureBuf_721;
         Mult_Buf[35].Weight_n = Wgt_7_721;
         Mult_Buf[36].Feature_n = FeatureBuf_722;
         Mult_Buf[36].Weight_n = Wgt_7_722;
         Mult_Buf[37].Feature_n = FeatureBuf_723;
         Mult_Buf[37].Weight_n = Wgt_7_723;
         Mult_Buf[38].Feature_n = FeatureBuf_724;
         Mult_Buf[38].Weight_n = Wgt_7_724;
         Mult_Buf[39].Feature_n = FeatureBuf_725;
         Mult_Buf[39].Weight_n = Wgt_7_725;
         Mult_Buf[40].Feature_n = FeatureBuf_726;
         Mult_Buf[40].Weight_n = Wgt_7_726;
         Mult_Buf[41].Feature_n = FeatureBuf_727;
         Mult_Buf[41].Weight_n = Wgt_7_727;
         Mult_Buf[42].Feature_n = FeatureBuf_728;
         Mult_Buf[42].Weight_n = Wgt_7_728;
         Mult_Buf[43].Feature_n = FeatureBuf_729;
         Mult_Buf[43].Weight_n = Wgt_7_729;
         Mult_Buf[44].Feature_n = FeatureBuf_730;
         Mult_Buf[44].Weight_n = Wgt_7_730;
         Mult_Buf[45].Feature_n = FeatureBuf_731;
         Mult_Buf[45].Weight_n = Wgt_7_731;
         Mult_Buf[46].Feature_n = FeatureBuf_732;
         Mult_Buf[46].Weight_n = Wgt_7_732;
         Mult_Buf[47].Feature_n = FeatureBuf_733;
         Mult_Buf[47].Weight_n = Wgt_7_733;
         Mult_Buf[48].Feature_n = FeatureBuf_734;
         Mult_Buf[48].Weight_n = Wgt_7_734;
         Mult_Buf[49].Feature_n = FeatureBuf_735;
         Mult_Buf[49].Weight_n = Wgt_7_735;
         Mult_Buf[50].Feature_n = FeatureBuf_736;
         Mult_Buf[50].Weight_n = Wgt_7_736;
         Mult_Buf[51].Feature_n = FeatureBuf_737;
         Mult_Buf[51].Weight_n = Wgt_7_737;
         Mult_Buf[52].Feature_n = FeatureBuf_738;
         Mult_Buf[52].Weight_n = Wgt_7_738;
         Mult_Buf[53].Feature_n = FeatureBuf_739;
         Mult_Buf[53].Weight_n = Wgt_7_739;
         Mult_Buf[54].Feature_n = FeatureBuf_740;
         Mult_Buf[54].Weight_n = Wgt_7_740;
         Mult_Buf[55].Feature_n = FeatureBuf_741;
         Mult_Buf[55].Weight_n = Wgt_7_741;
         Mult_Buf[56].Feature_n = FeatureBuf_742;
         Mult_Buf[56].Weight_n = Wgt_7_742;
         Mult_Buf[57].Feature_n = FeatureBuf_743;
         Mult_Buf[57].Weight_n = Wgt_7_743;
         Mult_Buf[58].Feature_n = FeatureBuf_744;
         Mult_Buf[58].Weight_n = Wgt_7_744;
         Mult_Buf[59].Feature_n = FeatureBuf_745;
         Mult_Buf[59].Weight_n = Wgt_7_745;
         Mult_Buf[60].Feature_n = FeatureBuf_746;
         Mult_Buf[60].Weight_n = Wgt_7_746;
         Mult_Buf[61].Feature_n = FeatureBuf_747;
         Mult_Buf[61].Weight_n = Wgt_7_747;
         Mult_Buf[62].Feature_n = FeatureBuf_748;
         Mult_Buf[62].Weight_n = Wgt_7_748;
         Mult_Buf[63].Feature_n = FeatureBuf_749;
         Mult_Buf[63].Weight_n = Wgt_7_749;
         Mult_Buf[64].Feature_n = FeatureBuf_750;
         Mult_Buf[64].Weight_n = Wgt_7_750;
         Mult_Buf[65].Feature_n = FeatureBuf_751;
         Mult_Buf[65].Weight_n = Wgt_7_751;
         Mult_Buf[66].Feature_n = FeatureBuf_752;
         Mult_Buf[66].Weight_n = Wgt_7_752;
         Mult_Buf[67].Feature_n = FeatureBuf_753;
         Mult_Buf[67].Weight_n = Wgt_7_753;
         Mult_Buf[68].Feature_n = FeatureBuf_754;
         Mult_Buf[68].Weight_n = Wgt_7_754;
         Mult_Buf[69].Feature_n = FeatureBuf_755;
         Mult_Buf[69].Weight_n = Wgt_7_755;
         Mult_Buf[70].Feature_n = FeatureBuf_756;
         Mult_Buf[70].Weight_n = Wgt_7_756;
         Mult_Buf[71].Feature_n = FeatureBuf_757;
         Mult_Buf[71].Weight_n = Wgt_7_757;
         Mult_Buf[72].Feature_n = FeatureBuf_758;
         Mult_Buf[72].Weight_n = Wgt_7_758;
         Mult_Buf[73].Feature_n = FeatureBuf_759;
         Mult_Buf[73].Weight_n = Wgt_7_759;
         Mult_Buf[74].Feature_n = FeatureBuf_760;
         Mult_Buf[74].Weight_n = Wgt_7_760;
         Mult_Buf[75].Feature_n = FeatureBuf_761;
         Mult_Buf[75].Weight_n = Wgt_7_761;
         Mult_Buf[76].Feature_n = FeatureBuf_762;
         Mult_Buf[76].Weight_n = Wgt_7_762;
         Mult_Buf[77].Feature_n = FeatureBuf_763;
         Mult_Buf[77].Weight_n = Wgt_7_763;
         Mult_Buf[78].Feature_n = FeatureBuf_764;
         Mult_Buf[78].Weight_n = Wgt_7_764;
         Mult_Buf[79].Feature_n = FeatureBuf_765;
         Mult_Buf[79].Weight_n = Wgt_7_765;
         Mult_Buf[80].Feature_n = FeatureBuf_766;
         Mult_Buf[80].Weight_n = Wgt_7_766;
         Mult_Buf[81].Feature_n = FeatureBuf_767;
         Mult_Buf[81].Weight_n = Wgt_7_767;
         Mult_Buf[82].Feature_n = FeatureBuf_768;
         Mult_Buf[82].Weight_n = Wgt_7_768;
         Mult_Buf[83].Feature_n = FeatureBuf_769;
         Mult_Buf[83].Weight_n = Wgt_7_769;
         Mult_Buf[84].Feature_n = FeatureBuf_770;
         Mult_Buf[84].Weight_n = Wgt_7_770;
         Mult_Buf[85].Feature_n = FeatureBuf_771;
         Mult_Buf[85].Weight_n = Wgt_7_771;
         Mult_Buf[86].Feature_n = FeatureBuf_772;
         Mult_Buf[86].Weight_n = Wgt_7_772;
         Mult_Buf[87].Feature_n = FeatureBuf_773;
         Mult_Buf[87].Weight_n = Wgt_7_773;
         Mult_Buf[88].Feature_n = FeatureBuf_774;
         Mult_Buf[88].Weight_n = Wgt_7_774;
         Mult_Buf[89].Feature_n = FeatureBuf_775;
         Mult_Buf[89].Weight_n = Wgt_7_775;
         Mult_Buf[90].Feature_n = FeatureBuf_776;
         Mult_Buf[90].Weight_n = Wgt_7_776;
         Mult_Buf[91].Feature_n = FeatureBuf_777;
         Mult_Buf[91].Weight_n = Wgt_7_777;
         Mult_Buf[92].Feature_n = FeatureBuf_778;
         Mult_Buf[92].Weight_n = Wgt_7_778;
         Mult_Buf[93].Feature_n = FeatureBuf_779;
         Mult_Buf[93].Weight_n = Wgt_7_779;
         Mult_Buf[94].Feature_n = FeatureBuf_780;
         Mult_Buf[94].Weight_n = Wgt_7_780;
         Mult_Buf[95].Feature_n = FeatureBuf_781;
         Mult_Buf[95].Weight_n = Wgt_7_781;
         Mult_Buf[96].Feature_n = FeatureBuf_782;
         Mult_Buf[96].Weight_n = Wgt_7_782;
         Mult_Buf[97].Feature_n = FeatureBuf_783;
         Mult_Buf[97].Weight_n = Wgt_7_783;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     //Collect Partial result form Adder
         Res_5_1_n = Part_Res;
     end
    66:begin
     nxt_state = 67;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_0;
         Mult_Buf[0].Weight_n = Wgt_8_0;
         Mult_Buf[1].Feature_n = FeatureBuf_1;
         Mult_Buf[1].Weight_n = Wgt_8_1;
         Mult_Buf[2].Feature_n = FeatureBuf_2;
         Mult_Buf[2].Weight_n = Wgt_8_2;
         Mult_Buf[3].Feature_n = FeatureBuf_3;
         Mult_Buf[3].Weight_n = Wgt_8_3;
         Mult_Buf[4].Feature_n = FeatureBuf_4;
         Mult_Buf[4].Weight_n = Wgt_8_4;
         Mult_Buf[5].Feature_n = FeatureBuf_5;
         Mult_Buf[5].Weight_n = Wgt_8_5;
         Mult_Buf[6].Feature_n = FeatureBuf_6;
         Mult_Buf[6].Weight_n = Wgt_8_6;
         Mult_Buf[7].Feature_n = FeatureBuf_7;
         Mult_Buf[7].Weight_n = Wgt_8_7;
         Mult_Buf[8].Feature_n = FeatureBuf_8;
         Mult_Buf[8].Weight_n = Wgt_8_8;
         Mult_Buf[9].Feature_n = FeatureBuf_9;
         Mult_Buf[9].Weight_n = Wgt_8_9;
         Mult_Buf[10].Feature_n = FeatureBuf_10;
         Mult_Buf[10].Weight_n = Wgt_8_10;
         Mult_Buf[11].Feature_n = FeatureBuf_11;
         Mult_Buf[11].Weight_n = Wgt_8_11;
         Mult_Buf[12].Feature_n = FeatureBuf_12;
         Mult_Buf[12].Weight_n = Wgt_8_12;
         Mult_Buf[13].Feature_n = FeatureBuf_13;
         Mult_Buf[13].Weight_n = Wgt_8_13;
         Mult_Buf[14].Feature_n = FeatureBuf_14;
         Mult_Buf[14].Weight_n = Wgt_8_14;
         Mult_Buf[15].Feature_n = FeatureBuf_15;
         Mult_Buf[15].Weight_n = Wgt_8_15;
         Mult_Buf[16].Feature_n = FeatureBuf_16;
         Mult_Buf[16].Weight_n = Wgt_8_16;
         Mult_Buf[17].Feature_n = FeatureBuf_17;
         Mult_Buf[17].Weight_n = Wgt_8_17;
         Mult_Buf[18].Feature_n = FeatureBuf_18;
         Mult_Buf[18].Weight_n = Wgt_8_18;
         Mult_Buf[19].Feature_n = FeatureBuf_19;
         Mult_Buf[19].Weight_n = Wgt_8_19;
         Mult_Buf[20].Feature_n = FeatureBuf_20;
         Mult_Buf[20].Weight_n = Wgt_8_20;
         Mult_Buf[21].Feature_n = FeatureBuf_21;
         Mult_Buf[21].Weight_n = Wgt_8_21;
         Mult_Buf[22].Feature_n = FeatureBuf_22;
         Mult_Buf[22].Weight_n = Wgt_8_22;
         Mult_Buf[23].Feature_n = FeatureBuf_23;
         Mult_Buf[23].Weight_n = Wgt_8_23;
         Mult_Buf[24].Feature_n = FeatureBuf_24;
         Mult_Buf[24].Weight_n = Wgt_8_24;
         Mult_Buf[25].Feature_n = FeatureBuf_25;
         Mult_Buf[25].Weight_n = Wgt_8_25;
         Mult_Buf[26].Feature_n = FeatureBuf_26;
         Mult_Buf[26].Weight_n = Wgt_8_26;
         Mult_Buf[27].Feature_n = FeatureBuf_27;
         Mult_Buf[27].Weight_n = Wgt_8_27;
         Mult_Buf[28].Feature_n = FeatureBuf_28;
         Mult_Buf[28].Weight_n = Wgt_8_28;
         Mult_Buf[29].Feature_n = FeatureBuf_29;
         Mult_Buf[29].Weight_n = Wgt_8_29;
         Mult_Buf[30].Feature_n = FeatureBuf_30;
         Mult_Buf[30].Weight_n = Wgt_8_30;
         Mult_Buf[31].Feature_n = FeatureBuf_31;
         Mult_Buf[31].Weight_n = Wgt_8_31;
         Mult_Buf[32].Feature_n = FeatureBuf_32;
         Mult_Buf[32].Weight_n = Wgt_8_32;
         Mult_Buf[33].Feature_n = FeatureBuf_33;
         Mult_Buf[33].Weight_n = Wgt_8_33;
         Mult_Buf[34].Feature_n = FeatureBuf_34;
         Mult_Buf[34].Weight_n = Wgt_8_34;
         Mult_Buf[35].Feature_n = FeatureBuf_35;
         Mult_Buf[35].Weight_n = Wgt_8_35;
         Mult_Buf[36].Feature_n = FeatureBuf_36;
         Mult_Buf[36].Weight_n = Wgt_8_36;
         Mult_Buf[37].Feature_n = FeatureBuf_37;
         Mult_Buf[37].Weight_n = Wgt_8_37;
         Mult_Buf[38].Feature_n = FeatureBuf_38;
         Mult_Buf[38].Weight_n = Wgt_8_38;
         Mult_Buf[39].Feature_n = FeatureBuf_39;
         Mult_Buf[39].Weight_n = Wgt_8_39;
         Mult_Buf[40].Feature_n = FeatureBuf_40;
         Mult_Buf[40].Weight_n = Wgt_8_40;
         Mult_Buf[41].Feature_n = FeatureBuf_41;
         Mult_Buf[41].Weight_n = Wgt_8_41;
         Mult_Buf[42].Feature_n = FeatureBuf_42;
         Mult_Buf[42].Weight_n = Wgt_8_42;
         Mult_Buf[43].Feature_n = FeatureBuf_43;
         Mult_Buf[43].Weight_n = Wgt_8_43;
         Mult_Buf[44].Feature_n = FeatureBuf_44;
         Mult_Buf[44].Weight_n = Wgt_8_44;
         Mult_Buf[45].Feature_n = FeatureBuf_45;
         Mult_Buf[45].Weight_n = Wgt_8_45;
         Mult_Buf[46].Feature_n = FeatureBuf_46;
         Mult_Buf[46].Weight_n = Wgt_8_46;
         Mult_Buf[47].Feature_n = FeatureBuf_47;
         Mult_Buf[47].Weight_n = Wgt_8_47;
         Mult_Buf[48].Feature_n = FeatureBuf_48;
         Mult_Buf[48].Weight_n = Wgt_8_48;
         Mult_Buf[49].Feature_n = FeatureBuf_49;
         Mult_Buf[49].Weight_n = Wgt_8_49;
         Mult_Buf[50].Feature_n = FeatureBuf_50;
         Mult_Buf[50].Weight_n = Wgt_8_50;
         Mult_Buf[51].Feature_n = FeatureBuf_51;
         Mult_Buf[51].Weight_n = Wgt_8_51;
         Mult_Buf[52].Feature_n = FeatureBuf_52;
         Mult_Buf[52].Weight_n = Wgt_8_52;
         Mult_Buf[53].Feature_n = FeatureBuf_53;
         Mult_Buf[53].Weight_n = Wgt_8_53;
         Mult_Buf[54].Feature_n = FeatureBuf_54;
         Mult_Buf[54].Weight_n = Wgt_8_54;
         Mult_Buf[55].Feature_n = FeatureBuf_55;
         Mult_Buf[55].Weight_n = Wgt_8_55;
         Mult_Buf[56].Feature_n = FeatureBuf_56;
         Mult_Buf[56].Weight_n = Wgt_8_56;
         Mult_Buf[57].Feature_n = FeatureBuf_57;
         Mult_Buf[57].Weight_n = Wgt_8_57;
         Mult_Buf[58].Feature_n = FeatureBuf_58;
         Mult_Buf[58].Weight_n = Wgt_8_58;
         Mult_Buf[59].Feature_n = FeatureBuf_59;
         Mult_Buf[59].Weight_n = Wgt_8_59;
         Mult_Buf[60].Feature_n = FeatureBuf_60;
         Mult_Buf[60].Weight_n = Wgt_8_60;
         Mult_Buf[61].Feature_n = FeatureBuf_61;
         Mult_Buf[61].Weight_n = Wgt_8_61;
         Mult_Buf[62].Feature_n = FeatureBuf_62;
         Mult_Buf[62].Weight_n = Wgt_8_62;
         Mult_Buf[63].Feature_n = FeatureBuf_63;
         Mult_Buf[63].Weight_n = Wgt_8_63;
         Mult_Buf[64].Feature_n = FeatureBuf_64;
         Mult_Buf[64].Weight_n = Wgt_8_64;
         Mult_Buf[65].Feature_n = FeatureBuf_65;
         Mult_Buf[65].Weight_n = Wgt_8_65;
         Mult_Buf[66].Feature_n = FeatureBuf_66;
         Mult_Buf[66].Weight_n = Wgt_8_66;
         Mult_Buf[67].Feature_n = FeatureBuf_67;
         Mult_Buf[67].Weight_n = Wgt_8_67;
         Mult_Buf[68].Feature_n = FeatureBuf_68;
         Mult_Buf[68].Weight_n = Wgt_8_68;
         Mult_Buf[69].Feature_n = FeatureBuf_69;
         Mult_Buf[69].Weight_n = Wgt_8_69;
         Mult_Buf[70].Feature_n = FeatureBuf_70;
         Mult_Buf[70].Weight_n = Wgt_8_70;
         Mult_Buf[71].Feature_n = FeatureBuf_71;
         Mult_Buf[71].Weight_n = Wgt_8_71;
         Mult_Buf[72].Feature_n = FeatureBuf_72;
         Mult_Buf[72].Weight_n = Wgt_8_72;
         Mult_Buf[73].Feature_n = FeatureBuf_73;
         Mult_Buf[73].Weight_n = Wgt_8_73;
         Mult_Buf[74].Feature_n = FeatureBuf_74;
         Mult_Buf[74].Weight_n = Wgt_8_74;
         Mult_Buf[75].Feature_n = FeatureBuf_75;
         Mult_Buf[75].Weight_n = Wgt_8_75;
         Mult_Buf[76].Feature_n = FeatureBuf_76;
         Mult_Buf[76].Weight_n = Wgt_8_76;
         Mult_Buf[77].Feature_n = FeatureBuf_77;
         Mult_Buf[77].Weight_n = Wgt_8_77;
         Mult_Buf[78].Feature_n = FeatureBuf_78;
         Mult_Buf[78].Weight_n = Wgt_8_78;
         Mult_Buf[79].Feature_n = FeatureBuf_79;
         Mult_Buf[79].Weight_n = Wgt_8_79;
         Mult_Buf[80].Feature_n = FeatureBuf_80;
         Mult_Buf[80].Weight_n = Wgt_8_80;
         Mult_Buf[81].Feature_n = FeatureBuf_81;
         Mult_Buf[81].Weight_n = Wgt_8_81;
         Mult_Buf[82].Feature_n = FeatureBuf_82;
         Mult_Buf[82].Weight_n = Wgt_8_82;
         Mult_Buf[83].Feature_n = FeatureBuf_83;
         Mult_Buf[83].Weight_n = Wgt_8_83;
         Mult_Buf[84].Feature_n = FeatureBuf_84;
         Mult_Buf[84].Weight_n = Wgt_8_84;
         Mult_Buf[85].Feature_n = FeatureBuf_85;
         Mult_Buf[85].Weight_n = Wgt_8_85;
         Mult_Buf[86].Feature_n = FeatureBuf_86;
         Mult_Buf[86].Weight_n = Wgt_8_86;
         Mult_Buf[87].Feature_n = FeatureBuf_87;
         Mult_Buf[87].Weight_n = Wgt_8_87;
         Mult_Buf[88].Feature_n = FeatureBuf_88;
         Mult_Buf[88].Weight_n = Wgt_8_88;
         Mult_Buf[89].Feature_n = FeatureBuf_89;
         Mult_Buf[89].Weight_n = Wgt_8_89;
         Mult_Buf[90].Feature_n = FeatureBuf_90;
         Mult_Buf[90].Weight_n = Wgt_8_90;
         Mult_Buf[91].Feature_n = FeatureBuf_91;
         Mult_Buf[91].Weight_n = Wgt_8_91;
         Mult_Buf[92].Feature_n = FeatureBuf_92;
         Mult_Buf[92].Weight_n = Wgt_8_92;
         Mult_Buf[93].Feature_n = FeatureBuf_93;
         Mult_Buf[93].Weight_n = Wgt_8_93;
         Mult_Buf[94].Feature_n = FeatureBuf_94;
         Mult_Buf[94].Weight_n = Wgt_8_94;
         Mult_Buf[95].Feature_n = FeatureBuf_95;
         Mult_Buf[95].Weight_n = Wgt_8_95;
         Mult_Buf[96].Feature_n = FeatureBuf_96;
         Mult_Buf[96].Weight_n = Wgt_8_96;
         Mult_Buf[97].Feature_n = FeatureBuf_97;
         Mult_Buf[97].Weight_n = Wgt_8_97;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     //Collect Partial result form Adder
         Res_5_2_n = Part_Res;
     end
    67:begin
     nxt_state = 68;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_98;
         Mult_Buf[0].Weight_n = Wgt_8_98;
         Mult_Buf[1].Feature_n = FeatureBuf_99;
         Mult_Buf[1].Weight_n = Wgt_8_99;
         Mult_Buf[2].Feature_n = FeatureBuf_100;
         Mult_Buf[2].Weight_n = Wgt_8_100;
         Mult_Buf[3].Feature_n = FeatureBuf_101;
         Mult_Buf[3].Weight_n = Wgt_8_101;
         Mult_Buf[4].Feature_n = FeatureBuf_102;
         Mult_Buf[4].Weight_n = Wgt_8_102;
         Mult_Buf[5].Feature_n = FeatureBuf_103;
         Mult_Buf[5].Weight_n = Wgt_8_103;
         Mult_Buf[6].Feature_n = FeatureBuf_104;
         Mult_Buf[6].Weight_n = Wgt_8_104;
         Mult_Buf[7].Feature_n = FeatureBuf_105;
         Mult_Buf[7].Weight_n = Wgt_8_105;
         Mult_Buf[8].Feature_n = FeatureBuf_106;
         Mult_Buf[8].Weight_n = Wgt_8_106;
         Mult_Buf[9].Feature_n = FeatureBuf_107;
         Mult_Buf[9].Weight_n = Wgt_8_107;
         Mult_Buf[10].Feature_n = FeatureBuf_108;
         Mult_Buf[10].Weight_n = Wgt_8_108;
         Mult_Buf[11].Feature_n = FeatureBuf_109;
         Mult_Buf[11].Weight_n = Wgt_8_109;
         Mult_Buf[12].Feature_n = FeatureBuf_110;
         Mult_Buf[12].Weight_n = Wgt_8_110;
         Mult_Buf[13].Feature_n = FeatureBuf_111;
         Mult_Buf[13].Weight_n = Wgt_8_111;
         Mult_Buf[14].Feature_n = FeatureBuf_112;
         Mult_Buf[14].Weight_n = Wgt_8_112;
         Mult_Buf[15].Feature_n = FeatureBuf_113;
         Mult_Buf[15].Weight_n = Wgt_8_113;
         Mult_Buf[16].Feature_n = FeatureBuf_114;
         Mult_Buf[16].Weight_n = Wgt_8_114;
         Mult_Buf[17].Feature_n = FeatureBuf_115;
         Mult_Buf[17].Weight_n = Wgt_8_115;
         Mult_Buf[18].Feature_n = FeatureBuf_116;
         Mult_Buf[18].Weight_n = Wgt_8_116;
         Mult_Buf[19].Feature_n = FeatureBuf_117;
         Mult_Buf[19].Weight_n = Wgt_8_117;
         Mult_Buf[20].Feature_n = FeatureBuf_118;
         Mult_Buf[20].Weight_n = Wgt_8_118;
         Mult_Buf[21].Feature_n = FeatureBuf_119;
         Mult_Buf[21].Weight_n = Wgt_8_119;
         Mult_Buf[22].Feature_n = FeatureBuf_120;
         Mult_Buf[22].Weight_n = Wgt_8_120;
         Mult_Buf[23].Feature_n = FeatureBuf_121;
         Mult_Buf[23].Weight_n = Wgt_8_121;
         Mult_Buf[24].Feature_n = FeatureBuf_122;
         Mult_Buf[24].Weight_n = Wgt_8_122;
         Mult_Buf[25].Feature_n = FeatureBuf_123;
         Mult_Buf[25].Weight_n = Wgt_8_123;
         Mult_Buf[26].Feature_n = FeatureBuf_124;
         Mult_Buf[26].Weight_n = Wgt_8_124;
         Mult_Buf[27].Feature_n = FeatureBuf_125;
         Mult_Buf[27].Weight_n = Wgt_8_125;
         Mult_Buf[28].Feature_n = FeatureBuf_126;
         Mult_Buf[28].Weight_n = Wgt_8_126;
         Mult_Buf[29].Feature_n = FeatureBuf_127;
         Mult_Buf[29].Weight_n = Wgt_8_127;
         Mult_Buf[30].Feature_n = FeatureBuf_128;
         Mult_Buf[30].Weight_n = Wgt_8_128;
         Mult_Buf[31].Feature_n = FeatureBuf_129;
         Mult_Buf[31].Weight_n = Wgt_8_129;
         Mult_Buf[32].Feature_n = FeatureBuf_130;
         Mult_Buf[32].Weight_n = Wgt_8_130;
         Mult_Buf[33].Feature_n = FeatureBuf_131;
         Mult_Buf[33].Weight_n = Wgt_8_131;
         Mult_Buf[34].Feature_n = FeatureBuf_132;
         Mult_Buf[34].Weight_n = Wgt_8_132;
         Mult_Buf[35].Feature_n = FeatureBuf_133;
         Mult_Buf[35].Weight_n = Wgt_8_133;
         Mult_Buf[36].Feature_n = FeatureBuf_134;
         Mult_Buf[36].Weight_n = Wgt_8_134;
         Mult_Buf[37].Feature_n = FeatureBuf_135;
         Mult_Buf[37].Weight_n = Wgt_8_135;
         Mult_Buf[38].Feature_n = FeatureBuf_136;
         Mult_Buf[38].Weight_n = Wgt_8_136;
         Mult_Buf[39].Feature_n = FeatureBuf_137;
         Mult_Buf[39].Weight_n = Wgt_8_137;
         Mult_Buf[40].Feature_n = FeatureBuf_138;
         Mult_Buf[40].Weight_n = Wgt_8_138;
         Mult_Buf[41].Feature_n = FeatureBuf_139;
         Mult_Buf[41].Weight_n = Wgt_8_139;
         Mult_Buf[42].Feature_n = FeatureBuf_140;
         Mult_Buf[42].Weight_n = Wgt_8_140;
         Mult_Buf[43].Feature_n = FeatureBuf_141;
         Mult_Buf[43].Weight_n = Wgt_8_141;
         Mult_Buf[44].Feature_n = FeatureBuf_142;
         Mult_Buf[44].Weight_n = Wgt_8_142;
         Mult_Buf[45].Feature_n = FeatureBuf_143;
         Mult_Buf[45].Weight_n = Wgt_8_143;
         Mult_Buf[46].Feature_n = FeatureBuf_144;
         Mult_Buf[46].Weight_n = Wgt_8_144;
         Mult_Buf[47].Feature_n = FeatureBuf_145;
         Mult_Buf[47].Weight_n = Wgt_8_145;
         Mult_Buf[48].Feature_n = FeatureBuf_146;
         Mult_Buf[48].Weight_n = Wgt_8_146;
         Mult_Buf[49].Feature_n = FeatureBuf_147;
         Mult_Buf[49].Weight_n = Wgt_8_147;
         Mult_Buf[50].Feature_n = FeatureBuf_148;
         Mult_Buf[50].Weight_n = Wgt_8_148;
         Mult_Buf[51].Feature_n = FeatureBuf_149;
         Mult_Buf[51].Weight_n = Wgt_8_149;
         Mult_Buf[52].Feature_n = FeatureBuf_150;
         Mult_Buf[52].Weight_n = Wgt_8_150;
         Mult_Buf[53].Feature_n = FeatureBuf_151;
         Mult_Buf[53].Weight_n = Wgt_8_151;
         Mult_Buf[54].Feature_n = FeatureBuf_152;
         Mult_Buf[54].Weight_n = Wgt_8_152;
         Mult_Buf[55].Feature_n = FeatureBuf_153;
         Mult_Buf[55].Weight_n = Wgt_8_153;
         Mult_Buf[56].Feature_n = FeatureBuf_154;
         Mult_Buf[56].Weight_n = Wgt_8_154;
         Mult_Buf[57].Feature_n = FeatureBuf_155;
         Mult_Buf[57].Weight_n = Wgt_8_155;
         Mult_Buf[58].Feature_n = FeatureBuf_156;
         Mult_Buf[58].Weight_n = Wgt_8_156;
         Mult_Buf[59].Feature_n = FeatureBuf_157;
         Mult_Buf[59].Weight_n = Wgt_8_157;
         Mult_Buf[60].Feature_n = FeatureBuf_158;
         Mult_Buf[60].Weight_n = Wgt_8_158;
         Mult_Buf[61].Feature_n = FeatureBuf_159;
         Mult_Buf[61].Weight_n = Wgt_8_159;
         Mult_Buf[62].Feature_n = FeatureBuf_160;
         Mult_Buf[62].Weight_n = Wgt_8_160;
         Mult_Buf[63].Feature_n = FeatureBuf_161;
         Mult_Buf[63].Weight_n = Wgt_8_161;
         Mult_Buf[64].Feature_n = FeatureBuf_162;
         Mult_Buf[64].Weight_n = Wgt_8_162;
         Mult_Buf[65].Feature_n = FeatureBuf_163;
         Mult_Buf[65].Weight_n = Wgt_8_163;
         Mult_Buf[66].Feature_n = FeatureBuf_164;
         Mult_Buf[66].Weight_n = Wgt_8_164;
         Mult_Buf[67].Feature_n = FeatureBuf_165;
         Mult_Buf[67].Weight_n = Wgt_8_165;
         Mult_Buf[68].Feature_n = FeatureBuf_166;
         Mult_Buf[68].Weight_n = Wgt_8_166;
         Mult_Buf[69].Feature_n = FeatureBuf_167;
         Mult_Buf[69].Weight_n = Wgt_8_167;
         Mult_Buf[70].Feature_n = FeatureBuf_168;
         Mult_Buf[70].Weight_n = Wgt_8_168;
         Mult_Buf[71].Feature_n = FeatureBuf_169;
         Mult_Buf[71].Weight_n = Wgt_8_169;
         Mult_Buf[72].Feature_n = FeatureBuf_170;
         Mult_Buf[72].Weight_n = Wgt_8_170;
         Mult_Buf[73].Feature_n = FeatureBuf_171;
         Mult_Buf[73].Weight_n = Wgt_8_171;
         Mult_Buf[74].Feature_n = FeatureBuf_172;
         Mult_Buf[74].Weight_n = Wgt_8_172;
         Mult_Buf[75].Feature_n = FeatureBuf_173;
         Mult_Buf[75].Weight_n = Wgt_8_173;
         Mult_Buf[76].Feature_n = FeatureBuf_174;
         Mult_Buf[76].Weight_n = Wgt_8_174;
         Mult_Buf[77].Feature_n = FeatureBuf_175;
         Mult_Buf[77].Weight_n = Wgt_8_175;
         Mult_Buf[78].Feature_n = FeatureBuf_176;
         Mult_Buf[78].Weight_n = Wgt_8_176;
         Mult_Buf[79].Feature_n = FeatureBuf_177;
         Mult_Buf[79].Weight_n = Wgt_8_177;
         Mult_Buf[80].Feature_n = FeatureBuf_178;
         Mult_Buf[80].Weight_n = Wgt_8_178;
         Mult_Buf[81].Feature_n = FeatureBuf_179;
         Mult_Buf[81].Weight_n = Wgt_8_179;
         Mult_Buf[82].Feature_n = FeatureBuf_180;
         Mult_Buf[82].Weight_n = Wgt_8_180;
         Mult_Buf[83].Feature_n = FeatureBuf_181;
         Mult_Buf[83].Weight_n = Wgt_8_181;
         Mult_Buf[84].Feature_n = FeatureBuf_182;
         Mult_Buf[84].Weight_n = Wgt_8_182;
         Mult_Buf[85].Feature_n = FeatureBuf_183;
         Mult_Buf[85].Weight_n = Wgt_8_183;
         Mult_Buf[86].Feature_n = FeatureBuf_184;
         Mult_Buf[86].Weight_n = Wgt_8_184;
         Mult_Buf[87].Feature_n = FeatureBuf_185;
         Mult_Buf[87].Weight_n = Wgt_8_185;
         Mult_Buf[88].Feature_n = FeatureBuf_186;
         Mult_Buf[88].Weight_n = Wgt_8_186;
         Mult_Buf[89].Feature_n = FeatureBuf_187;
         Mult_Buf[89].Weight_n = Wgt_8_187;
         Mult_Buf[90].Feature_n = FeatureBuf_188;
         Mult_Buf[90].Weight_n = Wgt_8_188;
         Mult_Buf[91].Feature_n = FeatureBuf_189;
         Mult_Buf[91].Weight_n = Wgt_8_189;
         Mult_Buf[92].Feature_n = FeatureBuf_190;
         Mult_Buf[92].Weight_n = Wgt_8_190;
         Mult_Buf[93].Feature_n = FeatureBuf_191;
         Mult_Buf[93].Weight_n = Wgt_8_191;
         Mult_Buf[94].Feature_n = FeatureBuf_192;
         Mult_Buf[94].Weight_n = Wgt_8_192;
         Mult_Buf[95].Feature_n = FeatureBuf_193;
         Mult_Buf[95].Weight_n = Wgt_8_193;
         Mult_Buf[96].Feature_n = FeatureBuf_194;
         Mult_Buf[96].Weight_n = Wgt_8_194;
         Mult_Buf[97].Feature_n = FeatureBuf_195;
         Mult_Buf[97].Weight_n = Wgt_8_195;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     //Collect Partial result form Adder
         Res_5_3_n = Part_Res;
     end
    68:begin
     nxt_state = 69;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_196;
         Mult_Buf[0].Weight_n = Wgt_8_196;
         Mult_Buf[1].Feature_n = FeatureBuf_197;
         Mult_Buf[1].Weight_n = Wgt_8_197;
         Mult_Buf[2].Feature_n = FeatureBuf_198;
         Mult_Buf[2].Weight_n = Wgt_8_198;
         Mult_Buf[3].Feature_n = FeatureBuf_199;
         Mult_Buf[3].Weight_n = Wgt_8_199;
         Mult_Buf[4].Feature_n = FeatureBuf_200;
         Mult_Buf[4].Weight_n = Wgt_8_200;
         Mult_Buf[5].Feature_n = FeatureBuf_201;
         Mult_Buf[5].Weight_n = Wgt_8_201;
         Mult_Buf[6].Feature_n = FeatureBuf_202;
         Mult_Buf[6].Weight_n = Wgt_8_202;
         Mult_Buf[7].Feature_n = FeatureBuf_203;
         Mult_Buf[7].Weight_n = Wgt_8_203;
         Mult_Buf[8].Feature_n = FeatureBuf_204;
         Mult_Buf[8].Weight_n = Wgt_8_204;
         Mult_Buf[9].Feature_n = FeatureBuf_205;
         Mult_Buf[9].Weight_n = Wgt_8_205;
         Mult_Buf[10].Feature_n = FeatureBuf_206;
         Mult_Buf[10].Weight_n = Wgt_8_206;
         Mult_Buf[11].Feature_n = FeatureBuf_207;
         Mult_Buf[11].Weight_n = Wgt_8_207;
         Mult_Buf[12].Feature_n = FeatureBuf_208;
         Mult_Buf[12].Weight_n = Wgt_8_208;
         Mult_Buf[13].Feature_n = FeatureBuf_209;
         Mult_Buf[13].Weight_n = Wgt_8_209;
         Mult_Buf[14].Feature_n = FeatureBuf_210;
         Mult_Buf[14].Weight_n = Wgt_8_210;
         Mult_Buf[15].Feature_n = FeatureBuf_211;
         Mult_Buf[15].Weight_n = Wgt_8_211;
         Mult_Buf[16].Feature_n = FeatureBuf_212;
         Mult_Buf[16].Weight_n = Wgt_8_212;
         Mult_Buf[17].Feature_n = FeatureBuf_213;
         Mult_Buf[17].Weight_n = Wgt_8_213;
         Mult_Buf[18].Feature_n = FeatureBuf_214;
         Mult_Buf[18].Weight_n = Wgt_8_214;
         Mult_Buf[19].Feature_n = FeatureBuf_215;
         Mult_Buf[19].Weight_n = Wgt_8_215;
         Mult_Buf[20].Feature_n = FeatureBuf_216;
         Mult_Buf[20].Weight_n = Wgt_8_216;
         Mult_Buf[21].Feature_n = FeatureBuf_217;
         Mult_Buf[21].Weight_n = Wgt_8_217;
         Mult_Buf[22].Feature_n = FeatureBuf_218;
         Mult_Buf[22].Weight_n = Wgt_8_218;
         Mult_Buf[23].Feature_n = FeatureBuf_219;
         Mult_Buf[23].Weight_n = Wgt_8_219;
         Mult_Buf[24].Feature_n = FeatureBuf_220;
         Mult_Buf[24].Weight_n = Wgt_8_220;
         Mult_Buf[25].Feature_n = FeatureBuf_221;
         Mult_Buf[25].Weight_n = Wgt_8_221;
         Mult_Buf[26].Feature_n = FeatureBuf_222;
         Mult_Buf[26].Weight_n = Wgt_8_222;
         Mult_Buf[27].Feature_n = FeatureBuf_223;
         Mult_Buf[27].Weight_n = Wgt_8_223;
         Mult_Buf[28].Feature_n = FeatureBuf_224;
         Mult_Buf[28].Weight_n = Wgt_8_224;
         Mult_Buf[29].Feature_n = FeatureBuf_225;
         Mult_Buf[29].Weight_n = Wgt_8_225;
         Mult_Buf[30].Feature_n = FeatureBuf_226;
         Mult_Buf[30].Weight_n = Wgt_8_226;
         Mult_Buf[31].Feature_n = FeatureBuf_227;
         Mult_Buf[31].Weight_n = Wgt_8_227;
         Mult_Buf[32].Feature_n = FeatureBuf_228;
         Mult_Buf[32].Weight_n = Wgt_8_228;
         Mult_Buf[33].Feature_n = FeatureBuf_229;
         Mult_Buf[33].Weight_n = Wgt_8_229;
         Mult_Buf[34].Feature_n = FeatureBuf_230;
         Mult_Buf[34].Weight_n = Wgt_8_230;
         Mult_Buf[35].Feature_n = FeatureBuf_231;
         Mult_Buf[35].Weight_n = Wgt_8_231;
         Mult_Buf[36].Feature_n = FeatureBuf_232;
         Mult_Buf[36].Weight_n = Wgt_8_232;
         Mult_Buf[37].Feature_n = FeatureBuf_233;
         Mult_Buf[37].Weight_n = Wgt_8_233;
         Mult_Buf[38].Feature_n = FeatureBuf_234;
         Mult_Buf[38].Weight_n = Wgt_8_234;
         Mult_Buf[39].Feature_n = FeatureBuf_235;
         Mult_Buf[39].Weight_n = Wgt_8_235;
         Mult_Buf[40].Feature_n = FeatureBuf_236;
         Mult_Buf[40].Weight_n = Wgt_8_236;
         Mult_Buf[41].Feature_n = FeatureBuf_237;
         Mult_Buf[41].Weight_n = Wgt_8_237;
         Mult_Buf[42].Feature_n = FeatureBuf_238;
         Mult_Buf[42].Weight_n = Wgt_8_238;
         Mult_Buf[43].Feature_n = FeatureBuf_239;
         Mult_Buf[43].Weight_n = Wgt_8_239;
         Mult_Buf[44].Feature_n = FeatureBuf_240;
         Mult_Buf[44].Weight_n = Wgt_8_240;
         Mult_Buf[45].Feature_n = FeatureBuf_241;
         Mult_Buf[45].Weight_n = Wgt_8_241;
         Mult_Buf[46].Feature_n = FeatureBuf_242;
         Mult_Buf[46].Weight_n = Wgt_8_242;
         Mult_Buf[47].Feature_n = FeatureBuf_243;
         Mult_Buf[47].Weight_n = Wgt_8_243;
         Mult_Buf[48].Feature_n = FeatureBuf_244;
         Mult_Buf[48].Weight_n = Wgt_8_244;
         Mult_Buf[49].Feature_n = FeatureBuf_245;
         Mult_Buf[49].Weight_n = Wgt_8_245;
         Mult_Buf[50].Feature_n = FeatureBuf_246;
         Mult_Buf[50].Weight_n = Wgt_8_246;
         Mult_Buf[51].Feature_n = FeatureBuf_247;
         Mult_Buf[51].Weight_n = Wgt_8_247;
         Mult_Buf[52].Feature_n = FeatureBuf_248;
         Mult_Buf[52].Weight_n = Wgt_8_248;
         Mult_Buf[53].Feature_n = FeatureBuf_249;
         Mult_Buf[53].Weight_n = Wgt_8_249;
         Mult_Buf[54].Feature_n = FeatureBuf_250;
         Mult_Buf[54].Weight_n = Wgt_8_250;
         Mult_Buf[55].Feature_n = FeatureBuf_251;
         Mult_Buf[55].Weight_n = Wgt_8_251;
         Mult_Buf[56].Feature_n = FeatureBuf_252;
         Mult_Buf[56].Weight_n = Wgt_8_252;
         Mult_Buf[57].Feature_n = FeatureBuf_253;
         Mult_Buf[57].Weight_n = Wgt_8_253;
         Mult_Buf[58].Feature_n = FeatureBuf_254;
         Mult_Buf[58].Weight_n = Wgt_8_254;
         Mult_Buf[59].Feature_n = FeatureBuf_255;
         Mult_Buf[59].Weight_n = Wgt_8_255;
         Mult_Buf[60].Feature_n = FeatureBuf_256;
         Mult_Buf[60].Weight_n = Wgt_8_256;
         Mult_Buf[61].Feature_n = FeatureBuf_257;
         Mult_Buf[61].Weight_n = Wgt_8_257;
         Mult_Buf[62].Feature_n = FeatureBuf_258;
         Mult_Buf[62].Weight_n = Wgt_8_258;
         Mult_Buf[63].Feature_n = FeatureBuf_259;
         Mult_Buf[63].Weight_n = Wgt_8_259;
         Mult_Buf[64].Feature_n = FeatureBuf_260;
         Mult_Buf[64].Weight_n = Wgt_8_260;
         Mult_Buf[65].Feature_n = FeatureBuf_261;
         Mult_Buf[65].Weight_n = Wgt_8_261;
         Mult_Buf[66].Feature_n = FeatureBuf_262;
         Mult_Buf[66].Weight_n = Wgt_8_262;
         Mult_Buf[67].Feature_n = FeatureBuf_263;
         Mult_Buf[67].Weight_n = Wgt_8_263;
         Mult_Buf[68].Feature_n = FeatureBuf_264;
         Mult_Buf[68].Weight_n = Wgt_8_264;
         Mult_Buf[69].Feature_n = FeatureBuf_265;
         Mult_Buf[69].Weight_n = Wgt_8_265;
         Mult_Buf[70].Feature_n = FeatureBuf_266;
         Mult_Buf[70].Weight_n = Wgt_8_266;
         Mult_Buf[71].Feature_n = FeatureBuf_267;
         Mult_Buf[71].Weight_n = Wgt_8_267;
         Mult_Buf[72].Feature_n = FeatureBuf_268;
         Mult_Buf[72].Weight_n = Wgt_8_268;
         Mult_Buf[73].Feature_n = FeatureBuf_269;
         Mult_Buf[73].Weight_n = Wgt_8_269;
         Mult_Buf[74].Feature_n = FeatureBuf_270;
         Mult_Buf[74].Weight_n = Wgt_8_270;
         Mult_Buf[75].Feature_n = FeatureBuf_271;
         Mult_Buf[75].Weight_n = Wgt_8_271;
         Mult_Buf[76].Feature_n = FeatureBuf_272;
         Mult_Buf[76].Weight_n = Wgt_8_272;
         Mult_Buf[77].Feature_n = FeatureBuf_273;
         Mult_Buf[77].Weight_n = Wgt_8_273;
         Mult_Buf[78].Feature_n = FeatureBuf_274;
         Mult_Buf[78].Weight_n = Wgt_8_274;
         Mult_Buf[79].Feature_n = FeatureBuf_275;
         Mult_Buf[79].Weight_n = Wgt_8_275;
         Mult_Buf[80].Feature_n = FeatureBuf_276;
         Mult_Buf[80].Weight_n = Wgt_8_276;
         Mult_Buf[81].Feature_n = FeatureBuf_277;
         Mult_Buf[81].Weight_n = Wgt_8_277;
         Mult_Buf[82].Feature_n = FeatureBuf_278;
         Mult_Buf[82].Weight_n = Wgt_8_278;
         Mult_Buf[83].Feature_n = FeatureBuf_279;
         Mult_Buf[83].Weight_n = Wgt_8_279;
         Mult_Buf[84].Feature_n = FeatureBuf_280;
         Mult_Buf[84].Weight_n = Wgt_8_280;
         Mult_Buf[85].Feature_n = FeatureBuf_281;
         Mult_Buf[85].Weight_n = Wgt_8_281;
         Mult_Buf[86].Feature_n = FeatureBuf_282;
         Mult_Buf[86].Weight_n = Wgt_8_282;
         Mult_Buf[87].Feature_n = FeatureBuf_283;
         Mult_Buf[87].Weight_n = Wgt_8_283;
         Mult_Buf[88].Feature_n = FeatureBuf_284;
         Mult_Buf[88].Weight_n = Wgt_8_284;
         Mult_Buf[89].Feature_n = FeatureBuf_285;
         Mult_Buf[89].Weight_n = Wgt_8_285;
         Mult_Buf[90].Feature_n = FeatureBuf_286;
         Mult_Buf[90].Weight_n = Wgt_8_286;
         Mult_Buf[91].Feature_n = FeatureBuf_287;
         Mult_Buf[91].Weight_n = Wgt_8_287;
         Mult_Buf[92].Feature_n = FeatureBuf_288;
         Mult_Buf[92].Weight_n = Wgt_8_288;
         Mult_Buf[93].Feature_n = FeatureBuf_289;
         Mult_Buf[93].Weight_n = Wgt_8_289;
         Mult_Buf[94].Feature_n = FeatureBuf_290;
         Mult_Buf[94].Weight_n = Wgt_8_290;
         Mult_Buf[95].Feature_n = FeatureBuf_291;
         Mult_Buf[95].Weight_n = Wgt_8_291;
         Mult_Buf[96].Feature_n = FeatureBuf_292;
         Mult_Buf[96].Weight_n = Wgt_8_292;
         Mult_Buf[97].Feature_n = FeatureBuf_293;
         Mult_Buf[97].Weight_n = Wgt_8_293;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     //Collect Partial result form Adder
         Res_5_4_n = Part_Res;
     end
    69:begin
     nxt_state = 70;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_294;
         Mult_Buf[0].Weight_n = Wgt_8_294;
         Mult_Buf[1].Feature_n = FeatureBuf_295;
         Mult_Buf[1].Weight_n = Wgt_8_295;
         Mult_Buf[2].Feature_n = FeatureBuf_296;
         Mult_Buf[2].Weight_n = Wgt_8_296;
         Mult_Buf[3].Feature_n = FeatureBuf_297;
         Mult_Buf[3].Weight_n = Wgt_8_297;
         Mult_Buf[4].Feature_n = FeatureBuf_298;
         Mult_Buf[4].Weight_n = Wgt_8_298;
         Mult_Buf[5].Feature_n = FeatureBuf_299;
         Mult_Buf[5].Weight_n = Wgt_8_299;
         Mult_Buf[6].Feature_n = FeatureBuf_300;
         Mult_Buf[6].Weight_n = Wgt_8_300;
         Mult_Buf[7].Feature_n = FeatureBuf_301;
         Mult_Buf[7].Weight_n = Wgt_8_301;
         Mult_Buf[8].Feature_n = FeatureBuf_302;
         Mult_Buf[8].Weight_n = Wgt_8_302;
         Mult_Buf[9].Feature_n = FeatureBuf_303;
         Mult_Buf[9].Weight_n = Wgt_8_303;
         Mult_Buf[10].Feature_n = FeatureBuf_304;
         Mult_Buf[10].Weight_n = Wgt_8_304;
         Mult_Buf[11].Feature_n = FeatureBuf_305;
         Mult_Buf[11].Weight_n = Wgt_8_305;
         Mult_Buf[12].Feature_n = FeatureBuf_306;
         Mult_Buf[12].Weight_n = Wgt_8_306;
         Mult_Buf[13].Feature_n = FeatureBuf_307;
         Mult_Buf[13].Weight_n = Wgt_8_307;
         Mult_Buf[14].Feature_n = FeatureBuf_308;
         Mult_Buf[14].Weight_n = Wgt_8_308;
         Mult_Buf[15].Feature_n = FeatureBuf_309;
         Mult_Buf[15].Weight_n = Wgt_8_309;
         Mult_Buf[16].Feature_n = FeatureBuf_310;
         Mult_Buf[16].Weight_n = Wgt_8_310;
         Mult_Buf[17].Feature_n = FeatureBuf_311;
         Mult_Buf[17].Weight_n = Wgt_8_311;
         Mult_Buf[18].Feature_n = FeatureBuf_312;
         Mult_Buf[18].Weight_n = Wgt_8_312;
         Mult_Buf[19].Feature_n = FeatureBuf_313;
         Mult_Buf[19].Weight_n = Wgt_8_313;
         Mult_Buf[20].Feature_n = FeatureBuf_314;
         Mult_Buf[20].Weight_n = Wgt_8_314;
         Mult_Buf[21].Feature_n = FeatureBuf_315;
         Mult_Buf[21].Weight_n = Wgt_8_315;
         Mult_Buf[22].Feature_n = FeatureBuf_316;
         Mult_Buf[22].Weight_n = Wgt_8_316;
         Mult_Buf[23].Feature_n = FeatureBuf_317;
         Mult_Buf[23].Weight_n = Wgt_8_317;
         Mult_Buf[24].Feature_n = FeatureBuf_318;
         Mult_Buf[24].Weight_n = Wgt_8_318;
         Mult_Buf[25].Feature_n = FeatureBuf_319;
         Mult_Buf[25].Weight_n = Wgt_8_319;
         Mult_Buf[26].Feature_n = FeatureBuf_320;
         Mult_Buf[26].Weight_n = Wgt_8_320;
         Mult_Buf[27].Feature_n = FeatureBuf_321;
         Mult_Buf[27].Weight_n = Wgt_8_321;
         Mult_Buf[28].Feature_n = FeatureBuf_322;
         Mult_Buf[28].Weight_n = Wgt_8_322;
         Mult_Buf[29].Feature_n = FeatureBuf_323;
         Mult_Buf[29].Weight_n = Wgt_8_323;
         Mult_Buf[30].Feature_n = FeatureBuf_324;
         Mult_Buf[30].Weight_n = Wgt_8_324;
         Mult_Buf[31].Feature_n = FeatureBuf_325;
         Mult_Buf[31].Weight_n = Wgt_8_325;
         Mult_Buf[32].Feature_n = FeatureBuf_326;
         Mult_Buf[32].Weight_n = Wgt_8_326;
         Mult_Buf[33].Feature_n = FeatureBuf_327;
         Mult_Buf[33].Weight_n = Wgt_8_327;
         Mult_Buf[34].Feature_n = FeatureBuf_328;
         Mult_Buf[34].Weight_n = Wgt_8_328;
         Mult_Buf[35].Feature_n = FeatureBuf_329;
         Mult_Buf[35].Weight_n = Wgt_8_329;
         Mult_Buf[36].Feature_n = FeatureBuf_330;
         Mult_Buf[36].Weight_n = Wgt_8_330;
         Mult_Buf[37].Feature_n = FeatureBuf_331;
         Mult_Buf[37].Weight_n = Wgt_8_331;
         Mult_Buf[38].Feature_n = FeatureBuf_332;
         Mult_Buf[38].Weight_n = Wgt_8_332;
         Mult_Buf[39].Feature_n = FeatureBuf_333;
         Mult_Buf[39].Weight_n = Wgt_8_333;
         Mult_Buf[40].Feature_n = FeatureBuf_334;
         Mult_Buf[40].Weight_n = Wgt_8_334;
         Mult_Buf[41].Feature_n = FeatureBuf_335;
         Mult_Buf[41].Weight_n = Wgt_8_335;
         Mult_Buf[42].Feature_n = FeatureBuf_336;
         Mult_Buf[42].Weight_n = Wgt_8_336;
         Mult_Buf[43].Feature_n = FeatureBuf_337;
         Mult_Buf[43].Weight_n = Wgt_8_337;
         Mult_Buf[44].Feature_n = FeatureBuf_338;
         Mult_Buf[44].Weight_n = Wgt_8_338;
         Mult_Buf[45].Feature_n = FeatureBuf_339;
         Mult_Buf[45].Weight_n = Wgt_8_339;
         Mult_Buf[46].Feature_n = FeatureBuf_340;
         Mult_Buf[46].Weight_n = Wgt_8_340;
         Mult_Buf[47].Feature_n = FeatureBuf_341;
         Mult_Buf[47].Weight_n = Wgt_8_341;
         Mult_Buf[48].Feature_n = FeatureBuf_342;
         Mult_Buf[48].Weight_n = Wgt_8_342;
         Mult_Buf[49].Feature_n = FeatureBuf_343;
         Mult_Buf[49].Weight_n = Wgt_8_343;
         Mult_Buf[50].Feature_n = FeatureBuf_344;
         Mult_Buf[50].Weight_n = Wgt_8_344;
         Mult_Buf[51].Feature_n = FeatureBuf_345;
         Mult_Buf[51].Weight_n = Wgt_8_345;
         Mult_Buf[52].Feature_n = FeatureBuf_346;
         Mult_Buf[52].Weight_n = Wgt_8_346;
         Mult_Buf[53].Feature_n = FeatureBuf_347;
         Mult_Buf[53].Weight_n = Wgt_8_347;
         Mult_Buf[54].Feature_n = FeatureBuf_348;
         Mult_Buf[54].Weight_n = Wgt_8_348;
         Mult_Buf[55].Feature_n = FeatureBuf_349;
         Mult_Buf[55].Weight_n = Wgt_8_349;
         Mult_Buf[56].Feature_n = FeatureBuf_350;
         Mult_Buf[56].Weight_n = Wgt_8_350;
         Mult_Buf[57].Feature_n = FeatureBuf_351;
         Mult_Buf[57].Weight_n = Wgt_8_351;
         Mult_Buf[58].Feature_n = FeatureBuf_352;
         Mult_Buf[58].Weight_n = Wgt_8_352;
         Mult_Buf[59].Feature_n = FeatureBuf_353;
         Mult_Buf[59].Weight_n = Wgt_8_353;
         Mult_Buf[60].Feature_n = FeatureBuf_354;
         Mult_Buf[60].Weight_n = Wgt_8_354;
         Mult_Buf[61].Feature_n = FeatureBuf_355;
         Mult_Buf[61].Weight_n = Wgt_8_355;
         Mult_Buf[62].Feature_n = FeatureBuf_356;
         Mult_Buf[62].Weight_n = Wgt_8_356;
         Mult_Buf[63].Feature_n = FeatureBuf_357;
         Mult_Buf[63].Weight_n = Wgt_8_357;
         Mult_Buf[64].Feature_n = FeatureBuf_358;
         Mult_Buf[64].Weight_n = Wgt_8_358;
         Mult_Buf[65].Feature_n = FeatureBuf_359;
         Mult_Buf[65].Weight_n = Wgt_8_359;
         Mult_Buf[66].Feature_n = FeatureBuf_360;
         Mult_Buf[66].Weight_n = Wgt_8_360;
         Mult_Buf[67].Feature_n = FeatureBuf_361;
         Mult_Buf[67].Weight_n = Wgt_8_361;
         Mult_Buf[68].Feature_n = FeatureBuf_362;
         Mult_Buf[68].Weight_n = Wgt_8_362;
         Mult_Buf[69].Feature_n = FeatureBuf_363;
         Mult_Buf[69].Weight_n = Wgt_8_363;
         Mult_Buf[70].Feature_n = FeatureBuf_364;
         Mult_Buf[70].Weight_n = Wgt_8_364;
         Mult_Buf[71].Feature_n = FeatureBuf_365;
         Mult_Buf[71].Weight_n = Wgt_8_365;
         Mult_Buf[72].Feature_n = FeatureBuf_366;
         Mult_Buf[72].Weight_n = Wgt_8_366;
         Mult_Buf[73].Feature_n = FeatureBuf_367;
         Mult_Buf[73].Weight_n = Wgt_8_367;
         Mult_Buf[74].Feature_n = FeatureBuf_368;
         Mult_Buf[74].Weight_n = Wgt_8_368;
         Mult_Buf[75].Feature_n = FeatureBuf_369;
         Mult_Buf[75].Weight_n = Wgt_8_369;
         Mult_Buf[76].Feature_n = FeatureBuf_370;
         Mult_Buf[76].Weight_n = Wgt_8_370;
         Mult_Buf[77].Feature_n = FeatureBuf_371;
         Mult_Buf[77].Weight_n = Wgt_8_371;
         Mult_Buf[78].Feature_n = FeatureBuf_372;
         Mult_Buf[78].Weight_n = Wgt_8_372;
         Mult_Buf[79].Feature_n = FeatureBuf_373;
         Mult_Buf[79].Weight_n = Wgt_8_373;
         Mult_Buf[80].Feature_n = FeatureBuf_374;
         Mult_Buf[80].Weight_n = Wgt_8_374;
         Mult_Buf[81].Feature_n = FeatureBuf_375;
         Mult_Buf[81].Weight_n = Wgt_8_375;
         Mult_Buf[82].Feature_n = FeatureBuf_376;
         Mult_Buf[82].Weight_n = Wgt_8_376;
         Mult_Buf[83].Feature_n = FeatureBuf_377;
         Mult_Buf[83].Weight_n = Wgt_8_377;
         Mult_Buf[84].Feature_n = FeatureBuf_378;
         Mult_Buf[84].Weight_n = Wgt_8_378;
         Mult_Buf[85].Feature_n = FeatureBuf_379;
         Mult_Buf[85].Weight_n = Wgt_8_379;
         Mult_Buf[86].Feature_n = FeatureBuf_380;
         Mult_Buf[86].Weight_n = Wgt_8_380;
         Mult_Buf[87].Feature_n = FeatureBuf_381;
         Mult_Buf[87].Weight_n = Wgt_8_381;
         Mult_Buf[88].Feature_n = FeatureBuf_382;
         Mult_Buf[88].Weight_n = Wgt_8_382;
         Mult_Buf[89].Feature_n = FeatureBuf_383;
         Mult_Buf[89].Weight_n = Wgt_8_383;
         Mult_Buf[90].Feature_n = FeatureBuf_384;
         Mult_Buf[90].Weight_n = Wgt_8_384;
         Mult_Buf[91].Feature_n = FeatureBuf_385;
         Mult_Buf[91].Weight_n = Wgt_8_385;
         Mult_Buf[92].Feature_n = FeatureBuf_386;
         Mult_Buf[92].Weight_n = Wgt_8_386;
         Mult_Buf[93].Feature_n = FeatureBuf_387;
         Mult_Buf[93].Weight_n = Wgt_8_387;
         Mult_Buf[94].Feature_n = FeatureBuf_388;
         Mult_Buf[94].Weight_n = Wgt_8_388;
         Mult_Buf[95].Feature_n = FeatureBuf_389;
         Mult_Buf[95].Weight_n = Wgt_8_389;
         Mult_Buf[96].Feature_n = FeatureBuf_390;
         Mult_Buf[96].Weight_n = Wgt_8_390;
         Mult_Buf[97].Feature_n = FeatureBuf_391;
         Mult_Buf[97].Weight_n = Wgt_8_391;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     //Collect Partial result form Adder
         Res_5_5_n = Part_Res;
     //Collect result from final Adder
         Res4_n = Final_Res;
     end
    70:begin
     nxt_state = 71;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_392;
         Mult_Buf[0].Weight_n = Wgt_8_392;
         Mult_Buf[1].Feature_n = FeatureBuf_393;
         Mult_Buf[1].Weight_n = Wgt_8_393;
         Mult_Buf[2].Feature_n = FeatureBuf_394;
         Mult_Buf[2].Weight_n = Wgt_8_394;
         Mult_Buf[3].Feature_n = FeatureBuf_395;
         Mult_Buf[3].Weight_n = Wgt_8_395;
         Mult_Buf[4].Feature_n = FeatureBuf_396;
         Mult_Buf[4].Weight_n = Wgt_8_396;
         Mult_Buf[5].Feature_n = FeatureBuf_397;
         Mult_Buf[5].Weight_n = Wgt_8_397;
         Mult_Buf[6].Feature_n = FeatureBuf_398;
         Mult_Buf[6].Weight_n = Wgt_8_398;
         Mult_Buf[7].Feature_n = FeatureBuf_399;
         Mult_Buf[7].Weight_n = Wgt_8_399;
         Mult_Buf[8].Feature_n = FeatureBuf_400;
         Mult_Buf[8].Weight_n = Wgt_8_400;
         Mult_Buf[9].Feature_n = FeatureBuf_401;
         Mult_Buf[9].Weight_n = Wgt_8_401;
         Mult_Buf[10].Feature_n = FeatureBuf_402;
         Mult_Buf[10].Weight_n = Wgt_8_402;
         Mult_Buf[11].Feature_n = FeatureBuf_403;
         Mult_Buf[11].Weight_n = Wgt_8_403;
         Mult_Buf[12].Feature_n = FeatureBuf_404;
         Mult_Buf[12].Weight_n = Wgt_8_404;
         Mult_Buf[13].Feature_n = FeatureBuf_405;
         Mult_Buf[13].Weight_n = Wgt_8_405;
         Mult_Buf[14].Feature_n = FeatureBuf_406;
         Mult_Buf[14].Weight_n = Wgt_8_406;
         Mult_Buf[15].Feature_n = FeatureBuf_407;
         Mult_Buf[15].Weight_n = Wgt_8_407;
         Mult_Buf[16].Feature_n = FeatureBuf_408;
         Mult_Buf[16].Weight_n = Wgt_8_408;
         Mult_Buf[17].Feature_n = FeatureBuf_409;
         Mult_Buf[17].Weight_n = Wgt_8_409;
         Mult_Buf[18].Feature_n = FeatureBuf_410;
         Mult_Buf[18].Weight_n = Wgt_8_410;
         Mult_Buf[19].Feature_n = FeatureBuf_411;
         Mult_Buf[19].Weight_n = Wgt_8_411;
         Mult_Buf[20].Feature_n = FeatureBuf_412;
         Mult_Buf[20].Weight_n = Wgt_8_412;
         Mult_Buf[21].Feature_n = FeatureBuf_413;
         Mult_Buf[21].Weight_n = Wgt_8_413;
         Mult_Buf[22].Feature_n = FeatureBuf_414;
         Mult_Buf[22].Weight_n = Wgt_8_414;
         Mult_Buf[23].Feature_n = FeatureBuf_415;
         Mult_Buf[23].Weight_n = Wgt_8_415;
         Mult_Buf[24].Feature_n = FeatureBuf_416;
         Mult_Buf[24].Weight_n = Wgt_8_416;
         Mult_Buf[25].Feature_n = FeatureBuf_417;
         Mult_Buf[25].Weight_n = Wgt_8_417;
         Mult_Buf[26].Feature_n = FeatureBuf_418;
         Mult_Buf[26].Weight_n = Wgt_8_418;
         Mult_Buf[27].Feature_n = FeatureBuf_419;
         Mult_Buf[27].Weight_n = Wgt_8_419;
         Mult_Buf[28].Feature_n = FeatureBuf_420;
         Mult_Buf[28].Weight_n = Wgt_8_420;
         Mult_Buf[29].Feature_n = FeatureBuf_421;
         Mult_Buf[29].Weight_n = Wgt_8_421;
         Mult_Buf[30].Feature_n = FeatureBuf_422;
         Mult_Buf[30].Weight_n = Wgt_8_422;
         Mult_Buf[31].Feature_n = FeatureBuf_423;
         Mult_Buf[31].Weight_n = Wgt_8_423;
         Mult_Buf[32].Feature_n = FeatureBuf_424;
         Mult_Buf[32].Weight_n = Wgt_8_424;
         Mult_Buf[33].Feature_n = FeatureBuf_425;
         Mult_Buf[33].Weight_n = Wgt_8_425;
         Mult_Buf[34].Feature_n = FeatureBuf_426;
         Mult_Buf[34].Weight_n = Wgt_8_426;
         Mult_Buf[35].Feature_n = FeatureBuf_427;
         Mult_Buf[35].Weight_n = Wgt_8_427;
         Mult_Buf[36].Feature_n = FeatureBuf_428;
         Mult_Buf[36].Weight_n = Wgt_8_428;
         Mult_Buf[37].Feature_n = FeatureBuf_429;
         Mult_Buf[37].Weight_n = Wgt_8_429;
         Mult_Buf[38].Feature_n = FeatureBuf_430;
         Mult_Buf[38].Weight_n = Wgt_8_430;
         Mult_Buf[39].Feature_n = FeatureBuf_431;
         Mult_Buf[39].Weight_n = Wgt_8_431;
         Mult_Buf[40].Feature_n = FeatureBuf_432;
         Mult_Buf[40].Weight_n = Wgt_8_432;
         Mult_Buf[41].Feature_n = FeatureBuf_433;
         Mult_Buf[41].Weight_n = Wgt_8_433;
         Mult_Buf[42].Feature_n = FeatureBuf_434;
         Mult_Buf[42].Weight_n = Wgt_8_434;
         Mult_Buf[43].Feature_n = FeatureBuf_435;
         Mult_Buf[43].Weight_n = Wgt_8_435;
         Mult_Buf[44].Feature_n = FeatureBuf_436;
         Mult_Buf[44].Weight_n = Wgt_8_436;
         Mult_Buf[45].Feature_n = FeatureBuf_437;
         Mult_Buf[45].Weight_n = Wgt_8_437;
         Mult_Buf[46].Feature_n = FeatureBuf_438;
         Mult_Buf[46].Weight_n = Wgt_8_438;
         Mult_Buf[47].Feature_n = FeatureBuf_439;
         Mult_Buf[47].Weight_n = Wgt_8_439;
         Mult_Buf[48].Feature_n = FeatureBuf_440;
         Mult_Buf[48].Weight_n = Wgt_8_440;
         Mult_Buf[49].Feature_n = FeatureBuf_441;
         Mult_Buf[49].Weight_n = Wgt_8_441;
         Mult_Buf[50].Feature_n = FeatureBuf_442;
         Mult_Buf[50].Weight_n = Wgt_8_442;
         Mult_Buf[51].Feature_n = FeatureBuf_443;
         Mult_Buf[51].Weight_n = Wgt_8_443;
         Mult_Buf[52].Feature_n = FeatureBuf_444;
         Mult_Buf[52].Weight_n = Wgt_8_444;
         Mult_Buf[53].Feature_n = FeatureBuf_445;
         Mult_Buf[53].Weight_n = Wgt_8_445;
         Mult_Buf[54].Feature_n = FeatureBuf_446;
         Mult_Buf[54].Weight_n = Wgt_8_446;
         Mult_Buf[55].Feature_n = FeatureBuf_447;
         Mult_Buf[55].Weight_n = Wgt_8_447;
         Mult_Buf[56].Feature_n = FeatureBuf_448;
         Mult_Buf[56].Weight_n = Wgt_8_448;
         Mult_Buf[57].Feature_n = FeatureBuf_449;
         Mult_Buf[57].Weight_n = Wgt_8_449;
         Mult_Buf[58].Feature_n = FeatureBuf_450;
         Mult_Buf[58].Weight_n = Wgt_8_450;
         Mult_Buf[59].Feature_n = FeatureBuf_451;
         Mult_Buf[59].Weight_n = Wgt_8_451;
         Mult_Buf[60].Feature_n = FeatureBuf_452;
         Mult_Buf[60].Weight_n = Wgt_8_452;
         Mult_Buf[61].Feature_n = FeatureBuf_453;
         Mult_Buf[61].Weight_n = Wgt_8_453;
         Mult_Buf[62].Feature_n = FeatureBuf_454;
         Mult_Buf[62].Weight_n = Wgt_8_454;
         Mult_Buf[63].Feature_n = FeatureBuf_455;
         Mult_Buf[63].Weight_n = Wgt_8_455;
         Mult_Buf[64].Feature_n = FeatureBuf_456;
         Mult_Buf[64].Weight_n = Wgt_8_456;
         Mult_Buf[65].Feature_n = FeatureBuf_457;
         Mult_Buf[65].Weight_n = Wgt_8_457;
         Mult_Buf[66].Feature_n = FeatureBuf_458;
         Mult_Buf[66].Weight_n = Wgt_8_458;
         Mult_Buf[67].Feature_n = FeatureBuf_459;
         Mult_Buf[67].Weight_n = Wgt_8_459;
         Mult_Buf[68].Feature_n = FeatureBuf_460;
         Mult_Buf[68].Weight_n = Wgt_8_460;
         Mult_Buf[69].Feature_n = FeatureBuf_461;
         Mult_Buf[69].Weight_n = Wgt_8_461;
         Mult_Buf[70].Feature_n = FeatureBuf_462;
         Mult_Buf[70].Weight_n = Wgt_8_462;
         Mult_Buf[71].Feature_n = FeatureBuf_463;
         Mult_Buf[71].Weight_n = Wgt_8_463;
         Mult_Buf[72].Feature_n = FeatureBuf_464;
         Mult_Buf[72].Weight_n = Wgt_8_464;
         Mult_Buf[73].Feature_n = FeatureBuf_465;
         Mult_Buf[73].Weight_n = Wgt_8_465;
         Mult_Buf[74].Feature_n = FeatureBuf_466;
         Mult_Buf[74].Weight_n = Wgt_8_466;
         Mult_Buf[75].Feature_n = FeatureBuf_467;
         Mult_Buf[75].Weight_n = Wgt_8_467;
         Mult_Buf[76].Feature_n = FeatureBuf_468;
         Mult_Buf[76].Weight_n = Wgt_8_468;
         Mult_Buf[77].Feature_n = FeatureBuf_469;
         Mult_Buf[77].Weight_n = Wgt_8_469;
         Mult_Buf[78].Feature_n = FeatureBuf_470;
         Mult_Buf[78].Weight_n = Wgt_8_470;
         Mult_Buf[79].Feature_n = FeatureBuf_471;
         Mult_Buf[79].Weight_n = Wgt_8_471;
         Mult_Buf[80].Feature_n = FeatureBuf_472;
         Mult_Buf[80].Weight_n = Wgt_8_472;
         Mult_Buf[81].Feature_n = FeatureBuf_473;
         Mult_Buf[81].Weight_n = Wgt_8_473;
         Mult_Buf[82].Feature_n = FeatureBuf_474;
         Mult_Buf[82].Weight_n = Wgt_8_474;
         Mult_Buf[83].Feature_n = FeatureBuf_475;
         Mult_Buf[83].Weight_n = Wgt_8_475;
         Mult_Buf[84].Feature_n = FeatureBuf_476;
         Mult_Buf[84].Weight_n = Wgt_8_476;
         Mult_Buf[85].Feature_n = FeatureBuf_477;
         Mult_Buf[85].Weight_n = Wgt_8_477;
         Mult_Buf[86].Feature_n = FeatureBuf_478;
         Mult_Buf[86].Weight_n = Wgt_8_478;
         Mult_Buf[87].Feature_n = FeatureBuf_479;
         Mult_Buf[87].Weight_n = Wgt_8_479;
         Mult_Buf[88].Feature_n = FeatureBuf_480;
         Mult_Buf[88].Weight_n = Wgt_8_480;
         Mult_Buf[89].Feature_n = FeatureBuf_481;
         Mult_Buf[89].Weight_n = Wgt_8_481;
         Mult_Buf[90].Feature_n = FeatureBuf_482;
         Mult_Buf[90].Weight_n = Wgt_8_482;
         Mult_Buf[91].Feature_n = FeatureBuf_483;
         Mult_Buf[91].Weight_n = Wgt_8_483;
         Mult_Buf[92].Feature_n = FeatureBuf_484;
         Mult_Buf[92].Weight_n = Wgt_8_484;
         Mult_Buf[93].Feature_n = FeatureBuf_485;
         Mult_Buf[93].Weight_n = Wgt_8_485;
         Mult_Buf[94].Feature_n = FeatureBuf_486;
         Mult_Buf[94].Weight_n = Wgt_8_486;
         Mult_Buf[95].Feature_n = FeatureBuf_487;
         Mult_Buf[95].Weight_n = Wgt_8_487;
         Mult_Buf[96].Feature_n = FeatureBuf_488;
         Mult_Buf[96].Weight_n = Wgt_8_488;
         Mult_Buf[97].Feature_n = FeatureBuf_489;
         Mult_Buf[97].Weight_n = Wgt_8_489;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     //Collect Partial result form Adder
         Res_5_6_n = Part_Res;
     end
    71:begin
     nxt_state = 72;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_490;
         Mult_Buf[0].Weight_n = Wgt_8_490;
         Mult_Buf[1].Feature_n = FeatureBuf_491;
         Mult_Buf[1].Weight_n = Wgt_8_491;
         Mult_Buf[2].Feature_n = FeatureBuf_492;
         Mult_Buf[2].Weight_n = Wgt_8_492;
         Mult_Buf[3].Feature_n = FeatureBuf_493;
         Mult_Buf[3].Weight_n = Wgt_8_493;
         Mult_Buf[4].Feature_n = FeatureBuf_494;
         Mult_Buf[4].Weight_n = Wgt_8_494;
         Mult_Buf[5].Feature_n = FeatureBuf_495;
         Mult_Buf[5].Weight_n = Wgt_8_495;
         Mult_Buf[6].Feature_n = FeatureBuf_496;
         Mult_Buf[6].Weight_n = Wgt_8_496;
         Mult_Buf[7].Feature_n = FeatureBuf_497;
         Mult_Buf[7].Weight_n = Wgt_8_497;
         Mult_Buf[8].Feature_n = FeatureBuf_498;
         Mult_Buf[8].Weight_n = Wgt_8_498;
         Mult_Buf[9].Feature_n = FeatureBuf_499;
         Mult_Buf[9].Weight_n = Wgt_8_499;
         Mult_Buf[10].Feature_n = FeatureBuf_500;
         Mult_Buf[10].Weight_n = Wgt_8_500;
         Mult_Buf[11].Feature_n = FeatureBuf_501;
         Mult_Buf[11].Weight_n = Wgt_8_501;
         Mult_Buf[12].Feature_n = FeatureBuf_502;
         Mult_Buf[12].Weight_n = Wgt_8_502;
         Mult_Buf[13].Feature_n = FeatureBuf_503;
         Mult_Buf[13].Weight_n = Wgt_8_503;
         Mult_Buf[14].Feature_n = FeatureBuf_504;
         Mult_Buf[14].Weight_n = Wgt_8_504;
         Mult_Buf[15].Feature_n = FeatureBuf_505;
         Mult_Buf[15].Weight_n = Wgt_8_505;
         Mult_Buf[16].Feature_n = FeatureBuf_506;
         Mult_Buf[16].Weight_n = Wgt_8_506;
         Mult_Buf[17].Feature_n = FeatureBuf_507;
         Mult_Buf[17].Weight_n = Wgt_8_507;
         Mult_Buf[18].Feature_n = FeatureBuf_508;
         Mult_Buf[18].Weight_n = Wgt_8_508;
         Mult_Buf[19].Feature_n = FeatureBuf_509;
         Mult_Buf[19].Weight_n = Wgt_8_509;
         Mult_Buf[20].Feature_n = FeatureBuf_510;
         Mult_Buf[20].Weight_n = Wgt_8_510;
         Mult_Buf[21].Feature_n = FeatureBuf_511;
         Mult_Buf[21].Weight_n = Wgt_8_511;
         Mult_Buf[22].Feature_n = FeatureBuf_512;
         Mult_Buf[22].Weight_n = Wgt_8_512;
         Mult_Buf[23].Feature_n = FeatureBuf_513;
         Mult_Buf[23].Weight_n = Wgt_8_513;
         Mult_Buf[24].Feature_n = FeatureBuf_514;
         Mult_Buf[24].Weight_n = Wgt_8_514;
         Mult_Buf[25].Feature_n = FeatureBuf_515;
         Mult_Buf[25].Weight_n = Wgt_8_515;
         Mult_Buf[26].Feature_n = FeatureBuf_516;
         Mult_Buf[26].Weight_n = Wgt_8_516;
         Mult_Buf[27].Feature_n = FeatureBuf_517;
         Mult_Buf[27].Weight_n = Wgt_8_517;
         Mult_Buf[28].Feature_n = FeatureBuf_518;
         Mult_Buf[28].Weight_n = Wgt_8_518;
         Mult_Buf[29].Feature_n = FeatureBuf_519;
         Mult_Buf[29].Weight_n = Wgt_8_519;
         Mult_Buf[30].Feature_n = FeatureBuf_520;
         Mult_Buf[30].Weight_n = Wgt_8_520;
         Mult_Buf[31].Feature_n = FeatureBuf_521;
         Mult_Buf[31].Weight_n = Wgt_8_521;
         Mult_Buf[32].Feature_n = FeatureBuf_522;
         Mult_Buf[32].Weight_n = Wgt_8_522;
         Mult_Buf[33].Feature_n = FeatureBuf_523;
         Mult_Buf[33].Weight_n = Wgt_8_523;
         Mult_Buf[34].Feature_n = FeatureBuf_524;
         Mult_Buf[34].Weight_n = Wgt_8_524;
         Mult_Buf[35].Feature_n = FeatureBuf_525;
         Mult_Buf[35].Weight_n = Wgt_8_525;
         Mult_Buf[36].Feature_n = FeatureBuf_526;
         Mult_Buf[36].Weight_n = Wgt_8_526;
         Mult_Buf[37].Feature_n = FeatureBuf_527;
         Mult_Buf[37].Weight_n = Wgt_8_527;
         Mult_Buf[38].Feature_n = FeatureBuf_528;
         Mult_Buf[38].Weight_n = Wgt_8_528;
         Mult_Buf[39].Feature_n = FeatureBuf_529;
         Mult_Buf[39].Weight_n = Wgt_8_529;
         Mult_Buf[40].Feature_n = FeatureBuf_530;
         Mult_Buf[40].Weight_n = Wgt_8_530;
         Mult_Buf[41].Feature_n = FeatureBuf_531;
         Mult_Buf[41].Weight_n = Wgt_8_531;
         Mult_Buf[42].Feature_n = FeatureBuf_532;
         Mult_Buf[42].Weight_n = Wgt_8_532;
         Mult_Buf[43].Feature_n = FeatureBuf_533;
         Mult_Buf[43].Weight_n = Wgt_8_533;
         Mult_Buf[44].Feature_n = FeatureBuf_534;
         Mult_Buf[44].Weight_n = Wgt_8_534;
         Mult_Buf[45].Feature_n = FeatureBuf_535;
         Mult_Buf[45].Weight_n = Wgt_8_535;
         Mult_Buf[46].Feature_n = FeatureBuf_536;
         Mult_Buf[46].Weight_n = Wgt_8_536;
         Mult_Buf[47].Feature_n = FeatureBuf_537;
         Mult_Buf[47].Weight_n = Wgt_8_537;
         Mult_Buf[48].Feature_n = FeatureBuf_538;
         Mult_Buf[48].Weight_n = Wgt_8_538;
         Mult_Buf[49].Feature_n = FeatureBuf_539;
         Mult_Buf[49].Weight_n = Wgt_8_539;
         Mult_Buf[50].Feature_n = FeatureBuf_540;
         Mult_Buf[50].Weight_n = Wgt_8_540;
         Mult_Buf[51].Feature_n = FeatureBuf_541;
         Mult_Buf[51].Weight_n = Wgt_8_541;
         Mult_Buf[52].Feature_n = FeatureBuf_542;
         Mult_Buf[52].Weight_n = Wgt_8_542;
         Mult_Buf[53].Feature_n = FeatureBuf_543;
         Mult_Buf[53].Weight_n = Wgt_8_543;
         Mult_Buf[54].Feature_n = FeatureBuf_544;
         Mult_Buf[54].Weight_n = Wgt_8_544;
         Mult_Buf[55].Feature_n = FeatureBuf_545;
         Mult_Buf[55].Weight_n = Wgt_8_545;
         Mult_Buf[56].Feature_n = FeatureBuf_546;
         Mult_Buf[56].Weight_n = Wgt_8_546;
         Mult_Buf[57].Feature_n = FeatureBuf_547;
         Mult_Buf[57].Weight_n = Wgt_8_547;
         Mult_Buf[58].Feature_n = FeatureBuf_548;
         Mult_Buf[58].Weight_n = Wgt_8_548;
         Mult_Buf[59].Feature_n = FeatureBuf_549;
         Mult_Buf[59].Weight_n = Wgt_8_549;
         Mult_Buf[60].Feature_n = FeatureBuf_550;
         Mult_Buf[60].Weight_n = Wgt_8_550;
         Mult_Buf[61].Feature_n = FeatureBuf_551;
         Mult_Buf[61].Weight_n = Wgt_8_551;
         Mult_Buf[62].Feature_n = FeatureBuf_552;
         Mult_Buf[62].Weight_n = Wgt_8_552;
         Mult_Buf[63].Feature_n = FeatureBuf_553;
         Mult_Buf[63].Weight_n = Wgt_8_553;
         Mult_Buf[64].Feature_n = FeatureBuf_554;
         Mult_Buf[64].Weight_n = Wgt_8_554;
         Mult_Buf[65].Feature_n = FeatureBuf_555;
         Mult_Buf[65].Weight_n = Wgt_8_555;
         Mult_Buf[66].Feature_n = FeatureBuf_556;
         Mult_Buf[66].Weight_n = Wgt_8_556;
         Mult_Buf[67].Feature_n = FeatureBuf_557;
         Mult_Buf[67].Weight_n = Wgt_8_557;
         Mult_Buf[68].Feature_n = FeatureBuf_558;
         Mult_Buf[68].Weight_n = Wgt_8_558;
         Mult_Buf[69].Feature_n = FeatureBuf_559;
         Mult_Buf[69].Weight_n = Wgt_8_559;
         Mult_Buf[70].Feature_n = FeatureBuf_560;
         Mult_Buf[70].Weight_n = Wgt_8_560;
         Mult_Buf[71].Feature_n = FeatureBuf_561;
         Mult_Buf[71].Weight_n = Wgt_8_561;
         Mult_Buf[72].Feature_n = FeatureBuf_562;
         Mult_Buf[72].Weight_n = Wgt_8_562;
         Mult_Buf[73].Feature_n = FeatureBuf_563;
         Mult_Buf[73].Weight_n = Wgt_8_563;
         Mult_Buf[74].Feature_n = FeatureBuf_564;
         Mult_Buf[74].Weight_n = Wgt_8_564;
         Mult_Buf[75].Feature_n = FeatureBuf_565;
         Mult_Buf[75].Weight_n = Wgt_8_565;
         Mult_Buf[76].Feature_n = FeatureBuf_566;
         Mult_Buf[76].Weight_n = Wgt_8_566;
         Mult_Buf[77].Feature_n = FeatureBuf_567;
         Mult_Buf[77].Weight_n = Wgt_8_567;
         Mult_Buf[78].Feature_n = FeatureBuf_568;
         Mult_Buf[78].Weight_n = Wgt_8_568;
         Mult_Buf[79].Feature_n = FeatureBuf_569;
         Mult_Buf[79].Weight_n = Wgt_8_569;
         Mult_Buf[80].Feature_n = FeatureBuf_570;
         Mult_Buf[80].Weight_n = Wgt_8_570;
         Mult_Buf[81].Feature_n = FeatureBuf_571;
         Mult_Buf[81].Weight_n = Wgt_8_571;
         Mult_Buf[82].Feature_n = FeatureBuf_572;
         Mult_Buf[82].Weight_n = Wgt_8_572;
         Mult_Buf[83].Feature_n = FeatureBuf_573;
         Mult_Buf[83].Weight_n = Wgt_8_573;
         Mult_Buf[84].Feature_n = FeatureBuf_574;
         Mult_Buf[84].Weight_n = Wgt_8_574;
         Mult_Buf[85].Feature_n = FeatureBuf_575;
         Mult_Buf[85].Weight_n = Wgt_8_575;
         Mult_Buf[86].Feature_n = FeatureBuf_576;
         Mult_Buf[86].Weight_n = Wgt_8_576;
         Mult_Buf[87].Feature_n = FeatureBuf_577;
         Mult_Buf[87].Weight_n = Wgt_8_577;
         Mult_Buf[88].Feature_n = FeatureBuf_578;
         Mult_Buf[88].Weight_n = Wgt_8_578;
         Mult_Buf[89].Feature_n = FeatureBuf_579;
         Mult_Buf[89].Weight_n = Wgt_8_579;
         Mult_Buf[90].Feature_n = FeatureBuf_580;
         Mult_Buf[90].Weight_n = Wgt_8_580;
         Mult_Buf[91].Feature_n = FeatureBuf_581;
         Mult_Buf[91].Weight_n = Wgt_8_581;
         Mult_Buf[92].Feature_n = FeatureBuf_582;
         Mult_Buf[92].Weight_n = Wgt_8_582;
         Mult_Buf[93].Feature_n = FeatureBuf_583;
         Mult_Buf[93].Weight_n = Wgt_8_583;
         Mult_Buf[94].Feature_n = FeatureBuf_584;
         Mult_Buf[94].Weight_n = Wgt_8_584;
         Mult_Buf[95].Feature_n = FeatureBuf_585;
         Mult_Buf[95].Weight_n = Wgt_8_585;
         Mult_Buf[96].Feature_n = FeatureBuf_586;
         Mult_Buf[96].Weight_n = Wgt_8_586;
         Mult_Buf[97].Feature_n = FeatureBuf_587;
         Mult_Buf[97].Weight_n = Wgt_8_587;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     //Collect Partial result form Adder
         Res_5_7_n = Part_Res;
     //Feed to final Adder
         A1 = Part_Res;
         A2 = Res_5_6_n;
         A3 = Res_5_5_n;
         A4 = Res_5_4_n;
         A5 = Res_5_3_n;
         A6 = Res_5_2_n;
         A7 = Res_5_1_n;
         A8 = Res_5_0_n;
     end
    72:begin
     nxt_state = 73;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_588;
         Mult_Buf[0].Weight_n = Wgt_8_588;
         Mult_Buf[1].Feature_n = FeatureBuf_589;
         Mult_Buf[1].Weight_n = Wgt_8_589;
         Mult_Buf[2].Feature_n = FeatureBuf_590;
         Mult_Buf[2].Weight_n = Wgt_8_590;
         Mult_Buf[3].Feature_n = FeatureBuf_591;
         Mult_Buf[3].Weight_n = Wgt_8_591;
         Mult_Buf[4].Feature_n = FeatureBuf_592;
         Mult_Buf[4].Weight_n = Wgt_8_592;
         Mult_Buf[5].Feature_n = FeatureBuf_593;
         Mult_Buf[5].Weight_n = Wgt_8_593;
         Mult_Buf[6].Feature_n = FeatureBuf_594;
         Mult_Buf[6].Weight_n = Wgt_8_594;
         Mult_Buf[7].Feature_n = FeatureBuf_595;
         Mult_Buf[7].Weight_n = Wgt_8_595;
         Mult_Buf[8].Feature_n = FeatureBuf_596;
         Mult_Buf[8].Weight_n = Wgt_8_596;
         Mult_Buf[9].Feature_n = FeatureBuf_597;
         Mult_Buf[9].Weight_n = Wgt_8_597;
         Mult_Buf[10].Feature_n = FeatureBuf_598;
         Mult_Buf[10].Weight_n = Wgt_8_598;
         Mult_Buf[11].Feature_n = FeatureBuf_599;
         Mult_Buf[11].Weight_n = Wgt_8_599;
         Mult_Buf[12].Feature_n = FeatureBuf_600;
         Mult_Buf[12].Weight_n = Wgt_8_600;
         Mult_Buf[13].Feature_n = FeatureBuf_601;
         Mult_Buf[13].Weight_n = Wgt_8_601;
         Mult_Buf[14].Feature_n = FeatureBuf_602;
         Mult_Buf[14].Weight_n = Wgt_8_602;
         Mult_Buf[15].Feature_n = FeatureBuf_603;
         Mult_Buf[15].Weight_n = Wgt_8_603;
         Mult_Buf[16].Feature_n = FeatureBuf_604;
         Mult_Buf[16].Weight_n = Wgt_8_604;
         Mult_Buf[17].Feature_n = FeatureBuf_605;
         Mult_Buf[17].Weight_n = Wgt_8_605;
         Mult_Buf[18].Feature_n = FeatureBuf_606;
         Mult_Buf[18].Weight_n = Wgt_8_606;
         Mult_Buf[19].Feature_n = FeatureBuf_607;
         Mult_Buf[19].Weight_n = Wgt_8_607;
         Mult_Buf[20].Feature_n = FeatureBuf_608;
         Mult_Buf[20].Weight_n = Wgt_8_608;
         Mult_Buf[21].Feature_n = FeatureBuf_609;
         Mult_Buf[21].Weight_n = Wgt_8_609;
         Mult_Buf[22].Feature_n = FeatureBuf_610;
         Mult_Buf[22].Weight_n = Wgt_8_610;
         Mult_Buf[23].Feature_n = FeatureBuf_611;
         Mult_Buf[23].Weight_n = Wgt_8_611;
         Mult_Buf[24].Feature_n = FeatureBuf_612;
         Mult_Buf[24].Weight_n = Wgt_8_612;
         Mult_Buf[25].Feature_n = FeatureBuf_613;
         Mult_Buf[25].Weight_n = Wgt_8_613;
         Mult_Buf[26].Feature_n = FeatureBuf_614;
         Mult_Buf[26].Weight_n = Wgt_8_614;
         Mult_Buf[27].Feature_n = FeatureBuf_615;
         Mult_Buf[27].Weight_n = Wgt_8_615;
         Mult_Buf[28].Feature_n = FeatureBuf_616;
         Mult_Buf[28].Weight_n = Wgt_8_616;
         Mult_Buf[29].Feature_n = FeatureBuf_617;
         Mult_Buf[29].Weight_n = Wgt_8_617;
         Mult_Buf[30].Feature_n = FeatureBuf_618;
         Mult_Buf[30].Weight_n = Wgt_8_618;
         Mult_Buf[31].Feature_n = FeatureBuf_619;
         Mult_Buf[31].Weight_n = Wgt_8_619;
         Mult_Buf[32].Feature_n = FeatureBuf_620;
         Mult_Buf[32].Weight_n = Wgt_8_620;
         Mult_Buf[33].Feature_n = FeatureBuf_621;
         Mult_Buf[33].Weight_n = Wgt_8_621;
         Mult_Buf[34].Feature_n = FeatureBuf_622;
         Mult_Buf[34].Weight_n = Wgt_8_622;
         Mult_Buf[35].Feature_n = FeatureBuf_623;
         Mult_Buf[35].Weight_n = Wgt_8_623;
         Mult_Buf[36].Feature_n = FeatureBuf_624;
         Mult_Buf[36].Weight_n = Wgt_8_624;
         Mult_Buf[37].Feature_n = FeatureBuf_625;
         Mult_Buf[37].Weight_n = Wgt_8_625;
         Mult_Buf[38].Feature_n = FeatureBuf_626;
         Mult_Buf[38].Weight_n = Wgt_8_626;
         Mult_Buf[39].Feature_n = FeatureBuf_627;
         Mult_Buf[39].Weight_n = Wgt_8_627;
         Mult_Buf[40].Feature_n = FeatureBuf_628;
         Mult_Buf[40].Weight_n = Wgt_8_628;
         Mult_Buf[41].Feature_n = FeatureBuf_629;
         Mult_Buf[41].Weight_n = Wgt_8_629;
         Mult_Buf[42].Feature_n = FeatureBuf_630;
         Mult_Buf[42].Weight_n = Wgt_8_630;
         Mult_Buf[43].Feature_n = FeatureBuf_631;
         Mult_Buf[43].Weight_n = Wgt_8_631;
         Mult_Buf[44].Feature_n = FeatureBuf_632;
         Mult_Buf[44].Weight_n = Wgt_8_632;
         Mult_Buf[45].Feature_n = FeatureBuf_633;
         Mult_Buf[45].Weight_n = Wgt_8_633;
         Mult_Buf[46].Feature_n = FeatureBuf_634;
         Mult_Buf[46].Weight_n = Wgt_8_634;
         Mult_Buf[47].Feature_n = FeatureBuf_635;
         Mult_Buf[47].Weight_n = Wgt_8_635;
         Mult_Buf[48].Feature_n = FeatureBuf_636;
         Mult_Buf[48].Weight_n = Wgt_8_636;
         Mult_Buf[49].Feature_n = FeatureBuf_637;
         Mult_Buf[49].Weight_n = Wgt_8_637;
         Mult_Buf[50].Feature_n = FeatureBuf_638;
         Mult_Buf[50].Weight_n = Wgt_8_638;
         Mult_Buf[51].Feature_n = FeatureBuf_639;
         Mult_Buf[51].Weight_n = Wgt_8_639;
         Mult_Buf[52].Feature_n = FeatureBuf_640;
         Mult_Buf[52].Weight_n = Wgt_8_640;
         Mult_Buf[53].Feature_n = FeatureBuf_641;
         Mult_Buf[53].Weight_n = Wgt_8_641;
         Mult_Buf[54].Feature_n = FeatureBuf_642;
         Mult_Buf[54].Weight_n = Wgt_8_642;
         Mult_Buf[55].Feature_n = FeatureBuf_643;
         Mult_Buf[55].Weight_n = Wgt_8_643;
         Mult_Buf[56].Feature_n = FeatureBuf_644;
         Mult_Buf[56].Weight_n = Wgt_8_644;
         Mult_Buf[57].Feature_n = FeatureBuf_645;
         Mult_Buf[57].Weight_n = Wgt_8_645;
         Mult_Buf[58].Feature_n = FeatureBuf_646;
         Mult_Buf[58].Weight_n = Wgt_8_646;
         Mult_Buf[59].Feature_n = FeatureBuf_647;
         Mult_Buf[59].Weight_n = Wgt_8_647;
         Mult_Buf[60].Feature_n = FeatureBuf_648;
         Mult_Buf[60].Weight_n = Wgt_8_648;
         Mult_Buf[61].Feature_n = FeatureBuf_649;
         Mult_Buf[61].Weight_n = Wgt_8_649;
         Mult_Buf[62].Feature_n = FeatureBuf_650;
         Mult_Buf[62].Weight_n = Wgt_8_650;
         Mult_Buf[63].Feature_n = FeatureBuf_651;
         Mult_Buf[63].Weight_n = Wgt_8_651;
         Mult_Buf[64].Feature_n = FeatureBuf_652;
         Mult_Buf[64].Weight_n = Wgt_8_652;
         Mult_Buf[65].Feature_n = FeatureBuf_653;
         Mult_Buf[65].Weight_n = Wgt_8_653;
         Mult_Buf[66].Feature_n = FeatureBuf_654;
         Mult_Buf[66].Weight_n = Wgt_8_654;
         Mult_Buf[67].Feature_n = FeatureBuf_655;
         Mult_Buf[67].Weight_n = Wgt_8_655;
         Mult_Buf[68].Feature_n = FeatureBuf_656;
         Mult_Buf[68].Weight_n = Wgt_8_656;
         Mult_Buf[69].Feature_n = FeatureBuf_657;
         Mult_Buf[69].Weight_n = Wgt_8_657;
         Mult_Buf[70].Feature_n = FeatureBuf_658;
         Mult_Buf[70].Weight_n = Wgt_8_658;
         Mult_Buf[71].Feature_n = FeatureBuf_659;
         Mult_Buf[71].Weight_n = Wgt_8_659;
         Mult_Buf[72].Feature_n = FeatureBuf_660;
         Mult_Buf[72].Weight_n = Wgt_8_660;
         Mult_Buf[73].Feature_n = FeatureBuf_661;
         Mult_Buf[73].Weight_n = Wgt_8_661;
         Mult_Buf[74].Feature_n = FeatureBuf_662;
         Mult_Buf[74].Weight_n = Wgt_8_662;
         Mult_Buf[75].Feature_n = FeatureBuf_663;
         Mult_Buf[75].Weight_n = Wgt_8_663;
         Mult_Buf[76].Feature_n = FeatureBuf_664;
         Mult_Buf[76].Weight_n = Wgt_8_664;
         Mult_Buf[77].Feature_n = FeatureBuf_665;
         Mult_Buf[77].Weight_n = Wgt_8_665;
         Mult_Buf[78].Feature_n = FeatureBuf_666;
         Mult_Buf[78].Weight_n = Wgt_8_666;
         Mult_Buf[79].Feature_n = FeatureBuf_667;
         Mult_Buf[79].Weight_n = Wgt_8_667;
         Mult_Buf[80].Feature_n = FeatureBuf_668;
         Mult_Buf[80].Weight_n = Wgt_8_668;
         Mult_Buf[81].Feature_n = FeatureBuf_669;
         Mult_Buf[81].Weight_n = Wgt_8_669;
         Mult_Buf[82].Feature_n = FeatureBuf_670;
         Mult_Buf[82].Weight_n = Wgt_8_670;
         Mult_Buf[83].Feature_n = FeatureBuf_671;
         Mult_Buf[83].Weight_n = Wgt_8_671;
         Mult_Buf[84].Feature_n = FeatureBuf_672;
         Mult_Buf[84].Weight_n = Wgt_8_672;
         Mult_Buf[85].Feature_n = FeatureBuf_673;
         Mult_Buf[85].Weight_n = Wgt_8_673;
         Mult_Buf[86].Feature_n = FeatureBuf_674;
         Mult_Buf[86].Weight_n = Wgt_8_674;
         Mult_Buf[87].Feature_n = FeatureBuf_675;
         Mult_Buf[87].Weight_n = Wgt_8_675;
         Mult_Buf[88].Feature_n = FeatureBuf_676;
         Mult_Buf[88].Weight_n = Wgt_8_676;
         Mult_Buf[89].Feature_n = FeatureBuf_677;
         Mult_Buf[89].Weight_n = Wgt_8_677;
         Mult_Buf[90].Feature_n = FeatureBuf_678;
         Mult_Buf[90].Weight_n = Wgt_8_678;
         Mult_Buf[91].Feature_n = FeatureBuf_679;
         Mult_Buf[91].Weight_n = Wgt_8_679;
         Mult_Buf[92].Feature_n = FeatureBuf_680;
         Mult_Buf[92].Weight_n = Wgt_8_680;
         Mult_Buf[93].Feature_n = FeatureBuf_681;
         Mult_Buf[93].Weight_n = Wgt_8_681;
         Mult_Buf[94].Feature_n = FeatureBuf_682;
         Mult_Buf[94].Weight_n = Wgt_8_682;
         Mult_Buf[95].Feature_n = FeatureBuf_683;
         Mult_Buf[95].Weight_n = Wgt_8_683;
         Mult_Buf[96].Feature_n = FeatureBuf_684;
         Mult_Buf[96].Weight_n = Wgt_8_684;
         Mult_Buf[97].Feature_n = FeatureBuf_685;
         Mult_Buf[97].Weight_n = Wgt_8_685;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     //Collect Partial result form Adder
         Res_6_0_n = Part_Res;
     end
    73:begin
     nxt_state = 74;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_686;
         Mult_Buf[0].Weight_n = Wgt_8_686;
         Mult_Buf[1].Feature_n = FeatureBuf_687;
         Mult_Buf[1].Weight_n = Wgt_8_687;
         Mult_Buf[2].Feature_n = FeatureBuf_688;
         Mult_Buf[2].Weight_n = Wgt_8_688;
         Mult_Buf[3].Feature_n = FeatureBuf_689;
         Mult_Buf[3].Weight_n = Wgt_8_689;
         Mult_Buf[4].Feature_n = FeatureBuf_690;
         Mult_Buf[4].Weight_n = Wgt_8_690;
         Mult_Buf[5].Feature_n = FeatureBuf_691;
         Mult_Buf[5].Weight_n = Wgt_8_691;
         Mult_Buf[6].Feature_n = FeatureBuf_692;
         Mult_Buf[6].Weight_n = Wgt_8_692;
         Mult_Buf[7].Feature_n = FeatureBuf_693;
         Mult_Buf[7].Weight_n = Wgt_8_693;
         Mult_Buf[8].Feature_n = FeatureBuf_694;
         Mult_Buf[8].Weight_n = Wgt_8_694;
         Mult_Buf[9].Feature_n = FeatureBuf_695;
         Mult_Buf[9].Weight_n = Wgt_8_695;
         Mult_Buf[10].Feature_n = FeatureBuf_696;
         Mult_Buf[10].Weight_n = Wgt_8_696;
         Mult_Buf[11].Feature_n = FeatureBuf_697;
         Mult_Buf[11].Weight_n = Wgt_8_697;
         Mult_Buf[12].Feature_n = FeatureBuf_698;
         Mult_Buf[12].Weight_n = Wgt_8_698;
         Mult_Buf[13].Feature_n = FeatureBuf_699;
         Mult_Buf[13].Weight_n = Wgt_8_699;
         Mult_Buf[14].Feature_n = FeatureBuf_700;
         Mult_Buf[14].Weight_n = Wgt_8_700;
         Mult_Buf[15].Feature_n = FeatureBuf_701;
         Mult_Buf[15].Weight_n = Wgt_8_701;
         Mult_Buf[16].Feature_n = FeatureBuf_702;
         Mult_Buf[16].Weight_n = Wgt_8_702;
         Mult_Buf[17].Feature_n = FeatureBuf_703;
         Mult_Buf[17].Weight_n = Wgt_8_703;
         Mult_Buf[18].Feature_n = FeatureBuf_704;
         Mult_Buf[18].Weight_n = Wgt_8_704;
         Mult_Buf[19].Feature_n = FeatureBuf_705;
         Mult_Buf[19].Weight_n = Wgt_8_705;
         Mult_Buf[20].Feature_n = FeatureBuf_706;
         Mult_Buf[20].Weight_n = Wgt_8_706;
         Mult_Buf[21].Feature_n = FeatureBuf_707;
         Mult_Buf[21].Weight_n = Wgt_8_707;
         Mult_Buf[22].Feature_n = FeatureBuf_708;
         Mult_Buf[22].Weight_n = Wgt_8_708;
         Mult_Buf[23].Feature_n = FeatureBuf_709;
         Mult_Buf[23].Weight_n = Wgt_8_709;
         Mult_Buf[24].Feature_n = FeatureBuf_710;
         Mult_Buf[24].Weight_n = Wgt_8_710;
         Mult_Buf[25].Feature_n = FeatureBuf_711;
         Mult_Buf[25].Weight_n = Wgt_8_711;
         Mult_Buf[26].Feature_n = FeatureBuf_712;
         Mult_Buf[26].Weight_n = Wgt_8_712;
         Mult_Buf[27].Feature_n = FeatureBuf_713;
         Mult_Buf[27].Weight_n = Wgt_8_713;
         Mult_Buf[28].Feature_n = FeatureBuf_714;
         Mult_Buf[28].Weight_n = Wgt_8_714;
         Mult_Buf[29].Feature_n = FeatureBuf_715;
         Mult_Buf[29].Weight_n = Wgt_8_715;
         Mult_Buf[30].Feature_n = FeatureBuf_716;
         Mult_Buf[30].Weight_n = Wgt_8_716;
         Mult_Buf[31].Feature_n = FeatureBuf_717;
         Mult_Buf[31].Weight_n = Wgt_8_717;
         Mult_Buf[32].Feature_n = FeatureBuf_718;
         Mult_Buf[32].Weight_n = Wgt_8_718;
         Mult_Buf[33].Feature_n = FeatureBuf_719;
         Mult_Buf[33].Weight_n = Wgt_8_719;
         Mult_Buf[34].Feature_n = FeatureBuf_720;
         Mult_Buf[34].Weight_n = Wgt_8_720;
         Mult_Buf[35].Feature_n = FeatureBuf_721;
         Mult_Buf[35].Weight_n = Wgt_8_721;
         Mult_Buf[36].Feature_n = FeatureBuf_722;
         Mult_Buf[36].Weight_n = Wgt_8_722;
         Mult_Buf[37].Feature_n = FeatureBuf_723;
         Mult_Buf[37].Weight_n = Wgt_8_723;
         Mult_Buf[38].Feature_n = FeatureBuf_724;
         Mult_Buf[38].Weight_n = Wgt_8_724;
         Mult_Buf[39].Feature_n = FeatureBuf_725;
         Mult_Buf[39].Weight_n = Wgt_8_725;
         Mult_Buf[40].Feature_n = FeatureBuf_726;
         Mult_Buf[40].Weight_n = Wgt_8_726;
         Mult_Buf[41].Feature_n = FeatureBuf_727;
         Mult_Buf[41].Weight_n = Wgt_8_727;
         Mult_Buf[42].Feature_n = FeatureBuf_728;
         Mult_Buf[42].Weight_n = Wgt_8_728;
         Mult_Buf[43].Feature_n = FeatureBuf_729;
         Mult_Buf[43].Weight_n = Wgt_8_729;
         Mult_Buf[44].Feature_n = FeatureBuf_730;
         Mult_Buf[44].Weight_n = Wgt_8_730;
         Mult_Buf[45].Feature_n = FeatureBuf_731;
         Mult_Buf[45].Weight_n = Wgt_8_731;
         Mult_Buf[46].Feature_n = FeatureBuf_732;
         Mult_Buf[46].Weight_n = Wgt_8_732;
         Mult_Buf[47].Feature_n = FeatureBuf_733;
         Mult_Buf[47].Weight_n = Wgt_8_733;
         Mult_Buf[48].Feature_n = FeatureBuf_734;
         Mult_Buf[48].Weight_n = Wgt_8_734;
         Mult_Buf[49].Feature_n = FeatureBuf_735;
         Mult_Buf[49].Weight_n = Wgt_8_735;
         Mult_Buf[50].Feature_n = FeatureBuf_736;
         Mult_Buf[50].Weight_n = Wgt_8_736;
         Mult_Buf[51].Feature_n = FeatureBuf_737;
         Mult_Buf[51].Weight_n = Wgt_8_737;
         Mult_Buf[52].Feature_n = FeatureBuf_738;
         Mult_Buf[52].Weight_n = Wgt_8_738;
         Mult_Buf[53].Feature_n = FeatureBuf_739;
         Mult_Buf[53].Weight_n = Wgt_8_739;
         Mult_Buf[54].Feature_n = FeatureBuf_740;
         Mult_Buf[54].Weight_n = Wgt_8_740;
         Mult_Buf[55].Feature_n = FeatureBuf_741;
         Mult_Buf[55].Weight_n = Wgt_8_741;
         Mult_Buf[56].Feature_n = FeatureBuf_742;
         Mult_Buf[56].Weight_n = Wgt_8_742;
         Mult_Buf[57].Feature_n = FeatureBuf_743;
         Mult_Buf[57].Weight_n = Wgt_8_743;
         Mult_Buf[58].Feature_n = FeatureBuf_744;
         Mult_Buf[58].Weight_n = Wgt_8_744;
         Mult_Buf[59].Feature_n = FeatureBuf_745;
         Mult_Buf[59].Weight_n = Wgt_8_745;
         Mult_Buf[60].Feature_n = FeatureBuf_746;
         Mult_Buf[60].Weight_n = Wgt_8_746;
         Mult_Buf[61].Feature_n = FeatureBuf_747;
         Mult_Buf[61].Weight_n = Wgt_8_747;
         Mult_Buf[62].Feature_n = FeatureBuf_748;
         Mult_Buf[62].Weight_n = Wgt_8_748;
         Mult_Buf[63].Feature_n = FeatureBuf_749;
         Mult_Buf[63].Weight_n = Wgt_8_749;
         Mult_Buf[64].Feature_n = FeatureBuf_750;
         Mult_Buf[64].Weight_n = Wgt_8_750;
         Mult_Buf[65].Feature_n = FeatureBuf_751;
         Mult_Buf[65].Weight_n = Wgt_8_751;
         Mult_Buf[66].Feature_n = FeatureBuf_752;
         Mult_Buf[66].Weight_n = Wgt_8_752;
         Mult_Buf[67].Feature_n = FeatureBuf_753;
         Mult_Buf[67].Weight_n = Wgt_8_753;
         Mult_Buf[68].Feature_n = FeatureBuf_754;
         Mult_Buf[68].Weight_n = Wgt_8_754;
         Mult_Buf[69].Feature_n = FeatureBuf_755;
         Mult_Buf[69].Weight_n = Wgt_8_755;
         Mult_Buf[70].Feature_n = FeatureBuf_756;
         Mult_Buf[70].Weight_n = Wgt_8_756;
         Mult_Buf[71].Feature_n = FeatureBuf_757;
         Mult_Buf[71].Weight_n = Wgt_8_757;
         Mult_Buf[72].Feature_n = FeatureBuf_758;
         Mult_Buf[72].Weight_n = Wgt_8_758;
         Mult_Buf[73].Feature_n = FeatureBuf_759;
         Mult_Buf[73].Weight_n = Wgt_8_759;
         Mult_Buf[74].Feature_n = FeatureBuf_760;
         Mult_Buf[74].Weight_n = Wgt_8_760;
         Mult_Buf[75].Feature_n = FeatureBuf_761;
         Mult_Buf[75].Weight_n = Wgt_8_761;
         Mult_Buf[76].Feature_n = FeatureBuf_762;
         Mult_Buf[76].Weight_n = Wgt_8_762;
         Mult_Buf[77].Feature_n = FeatureBuf_763;
         Mult_Buf[77].Weight_n = Wgt_8_763;
         Mult_Buf[78].Feature_n = FeatureBuf_764;
         Mult_Buf[78].Weight_n = Wgt_8_764;
         Mult_Buf[79].Feature_n = FeatureBuf_765;
         Mult_Buf[79].Weight_n = Wgt_8_765;
         Mult_Buf[80].Feature_n = FeatureBuf_766;
         Mult_Buf[80].Weight_n = Wgt_8_766;
         Mult_Buf[81].Feature_n = FeatureBuf_767;
         Mult_Buf[81].Weight_n = Wgt_8_767;
         Mult_Buf[82].Feature_n = FeatureBuf_768;
         Mult_Buf[82].Weight_n = Wgt_8_768;
         Mult_Buf[83].Feature_n = FeatureBuf_769;
         Mult_Buf[83].Weight_n = Wgt_8_769;
         Mult_Buf[84].Feature_n = FeatureBuf_770;
         Mult_Buf[84].Weight_n = Wgt_8_770;
         Mult_Buf[85].Feature_n = FeatureBuf_771;
         Mult_Buf[85].Weight_n = Wgt_8_771;
         Mult_Buf[86].Feature_n = FeatureBuf_772;
         Mult_Buf[86].Weight_n = Wgt_8_772;
         Mult_Buf[87].Feature_n = FeatureBuf_773;
         Mult_Buf[87].Weight_n = Wgt_8_773;
         Mult_Buf[88].Feature_n = FeatureBuf_774;
         Mult_Buf[88].Weight_n = Wgt_8_774;
         Mult_Buf[89].Feature_n = FeatureBuf_775;
         Mult_Buf[89].Weight_n = Wgt_8_775;
         Mult_Buf[90].Feature_n = FeatureBuf_776;
         Mult_Buf[90].Weight_n = Wgt_8_776;
         Mult_Buf[91].Feature_n = FeatureBuf_777;
         Mult_Buf[91].Weight_n = Wgt_8_777;
         Mult_Buf[92].Feature_n = FeatureBuf_778;
         Mult_Buf[92].Weight_n = Wgt_8_778;
         Mult_Buf[93].Feature_n = FeatureBuf_779;
         Mult_Buf[93].Weight_n = Wgt_8_779;
         Mult_Buf[94].Feature_n = FeatureBuf_780;
         Mult_Buf[94].Weight_n = Wgt_8_780;
         Mult_Buf[95].Feature_n = FeatureBuf_781;
         Mult_Buf[95].Weight_n = Wgt_8_781;
         Mult_Buf[96].Feature_n = FeatureBuf_782;
         Mult_Buf[96].Weight_n = Wgt_8_782;
         Mult_Buf[97].Feature_n = FeatureBuf_783;
         Mult_Buf[97].Weight_n = Wgt_8_783;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     //Collect Partial result form Adder
         Res_6_1_n = Part_Res;
     end
    74:begin
     nxt_state = 75;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_0;
         Mult_Buf[0].Weight_n = Wgt_9_0;
         Mult_Buf[1].Feature_n = FeatureBuf_1;
         Mult_Buf[1].Weight_n = Wgt_9_1;
         Mult_Buf[2].Feature_n = FeatureBuf_2;
         Mult_Buf[2].Weight_n = Wgt_9_2;
         Mult_Buf[3].Feature_n = FeatureBuf_3;
         Mult_Buf[3].Weight_n = Wgt_9_3;
         Mult_Buf[4].Feature_n = FeatureBuf_4;
         Mult_Buf[4].Weight_n = Wgt_9_4;
         Mult_Buf[5].Feature_n = FeatureBuf_5;
         Mult_Buf[5].Weight_n = Wgt_9_5;
         Mult_Buf[6].Feature_n = FeatureBuf_6;
         Mult_Buf[6].Weight_n = Wgt_9_6;
         Mult_Buf[7].Feature_n = FeatureBuf_7;
         Mult_Buf[7].Weight_n = Wgt_9_7;
         Mult_Buf[8].Feature_n = FeatureBuf_8;
         Mult_Buf[8].Weight_n = Wgt_9_8;
         Mult_Buf[9].Feature_n = FeatureBuf_9;
         Mult_Buf[9].Weight_n = Wgt_9_9;
         Mult_Buf[10].Feature_n = FeatureBuf_10;
         Mult_Buf[10].Weight_n = Wgt_9_10;
         Mult_Buf[11].Feature_n = FeatureBuf_11;
         Mult_Buf[11].Weight_n = Wgt_9_11;
         Mult_Buf[12].Feature_n = FeatureBuf_12;
         Mult_Buf[12].Weight_n = Wgt_9_12;
         Mult_Buf[13].Feature_n = FeatureBuf_13;
         Mult_Buf[13].Weight_n = Wgt_9_13;
         Mult_Buf[14].Feature_n = FeatureBuf_14;
         Mult_Buf[14].Weight_n = Wgt_9_14;
         Mult_Buf[15].Feature_n = FeatureBuf_15;
         Mult_Buf[15].Weight_n = Wgt_9_15;
         Mult_Buf[16].Feature_n = FeatureBuf_16;
         Mult_Buf[16].Weight_n = Wgt_9_16;
         Mult_Buf[17].Feature_n = FeatureBuf_17;
         Mult_Buf[17].Weight_n = Wgt_9_17;
         Mult_Buf[18].Feature_n = FeatureBuf_18;
         Mult_Buf[18].Weight_n = Wgt_9_18;
         Mult_Buf[19].Feature_n = FeatureBuf_19;
         Mult_Buf[19].Weight_n = Wgt_9_19;
         Mult_Buf[20].Feature_n = FeatureBuf_20;
         Mult_Buf[20].Weight_n = Wgt_9_20;
         Mult_Buf[21].Feature_n = FeatureBuf_21;
         Mult_Buf[21].Weight_n = Wgt_9_21;
         Mult_Buf[22].Feature_n = FeatureBuf_22;
         Mult_Buf[22].Weight_n = Wgt_9_22;
         Mult_Buf[23].Feature_n = FeatureBuf_23;
         Mult_Buf[23].Weight_n = Wgt_9_23;
         Mult_Buf[24].Feature_n = FeatureBuf_24;
         Mult_Buf[24].Weight_n = Wgt_9_24;
         Mult_Buf[25].Feature_n = FeatureBuf_25;
         Mult_Buf[25].Weight_n = Wgt_9_25;
         Mult_Buf[26].Feature_n = FeatureBuf_26;
         Mult_Buf[26].Weight_n = Wgt_9_26;
         Mult_Buf[27].Feature_n = FeatureBuf_27;
         Mult_Buf[27].Weight_n = Wgt_9_27;
         Mult_Buf[28].Feature_n = FeatureBuf_28;
         Mult_Buf[28].Weight_n = Wgt_9_28;
         Mult_Buf[29].Feature_n = FeatureBuf_29;
         Mult_Buf[29].Weight_n = Wgt_9_29;
         Mult_Buf[30].Feature_n = FeatureBuf_30;
         Mult_Buf[30].Weight_n = Wgt_9_30;
         Mult_Buf[31].Feature_n = FeatureBuf_31;
         Mult_Buf[31].Weight_n = Wgt_9_31;
         Mult_Buf[32].Feature_n = FeatureBuf_32;
         Mult_Buf[32].Weight_n = Wgt_9_32;
         Mult_Buf[33].Feature_n = FeatureBuf_33;
         Mult_Buf[33].Weight_n = Wgt_9_33;
         Mult_Buf[34].Feature_n = FeatureBuf_34;
         Mult_Buf[34].Weight_n = Wgt_9_34;
         Mult_Buf[35].Feature_n = FeatureBuf_35;
         Mult_Buf[35].Weight_n = Wgt_9_35;
         Mult_Buf[36].Feature_n = FeatureBuf_36;
         Mult_Buf[36].Weight_n = Wgt_9_36;
         Mult_Buf[37].Feature_n = FeatureBuf_37;
         Mult_Buf[37].Weight_n = Wgt_9_37;
         Mult_Buf[38].Feature_n = FeatureBuf_38;
         Mult_Buf[38].Weight_n = Wgt_9_38;
         Mult_Buf[39].Feature_n = FeatureBuf_39;
         Mult_Buf[39].Weight_n = Wgt_9_39;
         Mult_Buf[40].Feature_n = FeatureBuf_40;
         Mult_Buf[40].Weight_n = Wgt_9_40;
         Mult_Buf[41].Feature_n = FeatureBuf_41;
         Mult_Buf[41].Weight_n = Wgt_9_41;
         Mult_Buf[42].Feature_n = FeatureBuf_42;
         Mult_Buf[42].Weight_n = Wgt_9_42;
         Mult_Buf[43].Feature_n = FeatureBuf_43;
         Mult_Buf[43].Weight_n = Wgt_9_43;
         Mult_Buf[44].Feature_n = FeatureBuf_44;
         Mult_Buf[44].Weight_n = Wgt_9_44;
         Mult_Buf[45].Feature_n = FeatureBuf_45;
         Mult_Buf[45].Weight_n = Wgt_9_45;
         Mult_Buf[46].Feature_n = FeatureBuf_46;
         Mult_Buf[46].Weight_n = Wgt_9_46;
         Mult_Buf[47].Feature_n = FeatureBuf_47;
         Mult_Buf[47].Weight_n = Wgt_9_47;
         Mult_Buf[48].Feature_n = FeatureBuf_48;
         Mult_Buf[48].Weight_n = Wgt_9_48;
         Mult_Buf[49].Feature_n = FeatureBuf_49;
         Mult_Buf[49].Weight_n = Wgt_9_49;
         Mult_Buf[50].Feature_n = FeatureBuf_50;
         Mult_Buf[50].Weight_n = Wgt_9_50;
         Mult_Buf[51].Feature_n = FeatureBuf_51;
         Mult_Buf[51].Weight_n = Wgt_9_51;
         Mult_Buf[52].Feature_n = FeatureBuf_52;
         Mult_Buf[52].Weight_n = Wgt_9_52;
         Mult_Buf[53].Feature_n = FeatureBuf_53;
         Mult_Buf[53].Weight_n = Wgt_9_53;
         Mult_Buf[54].Feature_n = FeatureBuf_54;
         Mult_Buf[54].Weight_n = Wgt_9_54;
         Mult_Buf[55].Feature_n = FeatureBuf_55;
         Mult_Buf[55].Weight_n = Wgt_9_55;
         Mult_Buf[56].Feature_n = FeatureBuf_56;
         Mult_Buf[56].Weight_n = Wgt_9_56;
         Mult_Buf[57].Feature_n = FeatureBuf_57;
         Mult_Buf[57].Weight_n = Wgt_9_57;
         Mult_Buf[58].Feature_n = FeatureBuf_58;
         Mult_Buf[58].Weight_n = Wgt_9_58;
         Mult_Buf[59].Feature_n = FeatureBuf_59;
         Mult_Buf[59].Weight_n = Wgt_9_59;
         Mult_Buf[60].Feature_n = FeatureBuf_60;
         Mult_Buf[60].Weight_n = Wgt_9_60;
         Mult_Buf[61].Feature_n = FeatureBuf_61;
         Mult_Buf[61].Weight_n = Wgt_9_61;
         Mult_Buf[62].Feature_n = FeatureBuf_62;
         Mult_Buf[62].Weight_n = Wgt_9_62;
         Mult_Buf[63].Feature_n = FeatureBuf_63;
         Mult_Buf[63].Weight_n = Wgt_9_63;
         Mult_Buf[64].Feature_n = FeatureBuf_64;
         Mult_Buf[64].Weight_n = Wgt_9_64;
         Mult_Buf[65].Feature_n = FeatureBuf_65;
         Mult_Buf[65].Weight_n = Wgt_9_65;
         Mult_Buf[66].Feature_n = FeatureBuf_66;
         Mult_Buf[66].Weight_n = Wgt_9_66;
         Mult_Buf[67].Feature_n = FeatureBuf_67;
         Mult_Buf[67].Weight_n = Wgt_9_67;
         Mult_Buf[68].Feature_n = FeatureBuf_68;
         Mult_Buf[68].Weight_n = Wgt_9_68;
         Mult_Buf[69].Feature_n = FeatureBuf_69;
         Mult_Buf[69].Weight_n = Wgt_9_69;
         Mult_Buf[70].Feature_n = FeatureBuf_70;
         Mult_Buf[70].Weight_n = Wgt_9_70;
         Mult_Buf[71].Feature_n = FeatureBuf_71;
         Mult_Buf[71].Weight_n = Wgt_9_71;
         Mult_Buf[72].Feature_n = FeatureBuf_72;
         Mult_Buf[72].Weight_n = Wgt_9_72;
         Mult_Buf[73].Feature_n = FeatureBuf_73;
         Mult_Buf[73].Weight_n = Wgt_9_73;
         Mult_Buf[74].Feature_n = FeatureBuf_74;
         Mult_Buf[74].Weight_n = Wgt_9_74;
         Mult_Buf[75].Feature_n = FeatureBuf_75;
         Mult_Buf[75].Weight_n = Wgt_9_75;
         Mult_Buf[76].Feature_n = FeatureBuf_76;
         Mult_Buf[76].Weight_n = Wgt_9_76;
         Mult_Buf[77].Feature_n = FeatureBuf_77;
         Mult_Buf[77].Weight_n = Wgt_9_77;
         Mult_Buf[78].Feature_n = FeatureBuf_78;
         Mult_Buf[78].Weight_n = Wgt_9_78;
         Mult_Buf[79].Feature_n = FeatureBuf_79;
         Mult_Buf[79].Weight_n = Wgt_9_79;
         Mult_Buf[80].Feature_n = FeatureBuf_80;
         Mult_Buf[80].Weight_n = Wgt_9_80;
         Mult_Buf[81].Feature_n = FeatureBuf_81;
         Mult_Buf[81].Weight_n = Wgt_9_81;
         Mult_Buf[82].Feature_n = FeatureBuf_82;
         Mult_Buf[82].Weight_n = Wgt_9_82;
         Mult_Buf[83].Feature_n = FeatureBuf_83;
         Mult_Buf[83].Weight_n = Wgt_9_83;
         Mult_Buf[84].Feature_n = FeatureBuf_84;
         Mult_Buf[84].Weight_n = Wgt_9_84;
         Mult_Buf[85].Feature_n = FeatureBuf_85;
         Mult_Buf[85].Weight_n = Wgt_9_85;
         Mult_Buf[86].Feature_n = FeatureBuf_86;
         Mult_Buf[86].Weight_n = Wgt_9_86;
         Mult_Buf[87].Feature_n = FeatureBuf_87;
         Mult_Buf[87].Weight_n = Wgt_9_87;
         Mult_Buf[88].Feature_n = FeatureBuf_88;
         Mult_Buf[88].Weight_n = Wgt_9_88;
         Mult_Buf[89].Feature_n = FeatureBuf_89;
         Mult_Buf[89].Weight_n = Wgt_9_89;
         Mult_Buf[90].Feature_n = FeatureBuf_90;
         Mult_Buf[90].Weight_n = Wgt_9_90;
         Mult_Buf[91].Feature_n = FeatureBuf_91;
         Mult_Buf[91].Weight_n = Wgt_9_91;
         Mult_Buf[92].Feature_n = FeatureBuf_92;
         Mult_Buf[92].Weight_n = Wgt_9_92;
         Mult_Buf[93].Feature_n = FeatureBuf_93;
         Mult_Buf[93].Weight_n = Wgt_9_93;
         Mult_Buf[94].Feature_n = FeatureBuf_94;
         Mult_Buf[94].Weight_n = Wgt_9_94;
         Mult_Buf[95].Feature_n = FeatureBuf_95;
         Mult_Buf[95].Weight_n = Wgt_9_95;
         Mult_Buf[96].Feature_n = FeatureBuf_96;
         Mult_Buf[96].Weight_n = Wgt_9_96;
         Mult_Buf[97].Feature_n = FeatureBuf_97;
         Mult_Buf[97].Weight_n = Wgt_9_97;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     //Collect Partial result form Adder
         Res_6_2_n = Part_Res;
     end
    75:begin
     nxt_state = 76;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_98;
         Mult_Buf[0].Weight_n = Wgt_9_98;
         Mult_Buf[1].Feature_n = FeatureBuf_99;
         Mult_Buf[1].Weight_n = Wgt_9_99;
         Mult_Buf[2].Feature_n = FeatureBuf_100;
         Mult_Buf[2].Weight_n = Wgt_9_100;
         Mult_Buf[3].Feature_n = FeatureBuf_101;
         Mult_Buf[3].Weight_n = Wgt_9_101;
         Mult_Buf[4].Feature_n = FeatureBuf_102;
         Mult_Buf[4].Weight_n = Wgt_9_102;
         Mult_Buf[5].Feature_n = FeatureBuf_103;
         Mult_Buf[5].Weight_n = Wgt_9_103;
         Mult_Buf[6].Feature_n = FeatureBuf_104;
         Mult_Buf[6].Weight_n = Wgt_9_104;
         Mult_Buf[7].Feature_n = FeatureBuf_105;
         Mult_Buf[7].Weight_n = Wgt_9_105;
         Mult_Buf[8].Feature_n = FeatureBuf_106;
         Mult_Buf[8].Weight_n = Wgt_9_106;
         Mult_Buf[9].Feature_n = FeatureBuf_107;
         Mult_Buf[9].Weight_n = Wgt_9_107;
         Mult_Buf[10].Feature_n = FeatureBuf_108;
         Mult_Buf[10].Weight_n = Wgt_9_108;
         Mult_Buf[11].Feature_n = FeatureBuf_109;
         Mult_Buf[11].Weight_n = Wgt_9_109;
         Mult_Buf[12].Feature_n = FeatureBuf_110;
         Mult_Buf[12].Weight_n = Wgt_9_110;
         Mult_Buf[13].Feature_n = FeatureBuf_111;
         Mult_Buf[13].Weight_n = Wgt_9_111;
         Mult_Buf[14].Feature_n = FeatureBuf_112;
         Mult_Buf[14].Weight_n = Wgt_9_112;
         Mult_Buf[15].Feature_n = FeatureBuf_113;
         Mult_Buf[15].Weight_n = Wgt_9_113;
         Mult_Buf[16].Feature_n = FeatureBuf_114;
         Mult_Buf[16].Weight_n = Wgt_9_114;
         Mult_Buf[17].Feature_n = FeatureBuf_115;
         Mult_Buf[17].Weight_n = Wgt_9_115;
         Mult_Buf[18].Feature_n = FeatureBuf_116;
         Mult_Buf[18].Weight_n = Wgt_9_116;
         Mult_Buf[19].Feature_n = FeatureBuf_117;
         Mult_Buf[19].Weight_n = Wgt_9_117;
         Mult_Buf[20].Feature_n = FeatureBuf_118;
         Mult_Buf[20].Weight_n = Wgt_9_118;
         Mult_Buf[21].Feature_n = FeatureBuf_119;
         Mult_Buf[21].Weight_n = Wgt_9_119;
         Mult_Buf[22].Feature_n = FeatureBuf_120;
         Mult_Buf[22].Weight_n = Wgt_9_120;
         Mult_Buf[23].Feature_n = FeatureBuf_121;
         Mult_Buf[23].Weight_n = Wgt_9_121;
         Mult_Buf[24].Feature_n = FeatureBuf_122;
         Mult_Buf[24].Weight_n = Wgt_9_122;
         Mult_Buf[25].Feature_n = FeatureBuf_123;
         Mult_Buf[25].Weight_n = Wgt_9_123;
         Mult_Buf[26].Feature_n = FeatureBuf_124;
         Mult_Buf[26].Weight_n = Wgt_9_124;
         Mult_Buf[27].Feature_n = FeatureBuf_125;
         Mult_Buf[27].Weight_n = Wgt_9_125;
         Mult_Buf[28].Feature_n = FeatureBuf_126;
         Mult_Buf[28].Weight_n = Wgt_9_126;
         Mult_Buf[29].Feature_n = FeatureBuf_127;
         Mult_Buf[29].Weight_n = Wgt_9_127;
         Mult_Buf[30].Feature_n = FeatureBuf_128;
         Mult_Buf[30].Weight_n = Wgt_9_128;
         Mult_Buf[31].Feature_n = FeatureBuf_129;
         Mult_Buf[31].Weight_n = Wgt_9_129;
         Mult_Buf[32].Feature_n = FeatureBuf_130;
         Mult_Buf[32].Weight_n = Wgt_9_130;
         Mult_Buf[33].Feature_n = FeatureBuf_131;
         Mult_Buf[33].Weight_n = Wgt_9_131;
         Mult_Buf[34].Feature_n = FeatureBuf_132;
         Mult_Buf[34].Weight_n = Wgt_9_132;
         Mult_Buf[35].Feature_n = FeatureBuf_133;
         Mult_Buf[35].Weight_n = Wgt_9_133;
         Mult_Buf[36].Feature_n = FeatureBuf_134;
         Mult_Buf[36].Weight_n = Wgt_9_134;
         Mult_Buf[37].Feature_n = FeatureBuf_135;
         Mult_Buf[37].Weight_n = Wgt_9_135;
         Mult_Buf[38].Feature_n = FeatureBuf_136;
         Mult_Buf[38].Weight_n = Wgt_9_136;
         Mult_Buf[39].Feature_n = FeatureBuf_137;
         Mult_Buf[39].Weight_n = Wgt_9_137;
         Mult_Buf[40].Feature_n = FeatureBuf_138;
         Mult_Buf[40].Weight_n = Wgt_9_138;
         Mult_Buf[41].Feature_n = FeatureBuf_139;
         Mult_Buf[41].Weight_n = Wgt_9_139;
         Mult_Buf[42].Feature_n = FeatureBuf_140;
         Mult_Buf[42].Weight_n = Wgt_9_140;
         Mult_Buf[43].Feature_n = FeatureBuf_141;
         Mult_Buf[43].Weight_n = Wgt_9_141;
         Mult_Buf[44].Feature_n = FeatureBuf_142;
         Mult_Buf[44].Weight_n = Wgt_9_142;
         Mult_Buf[45].Feature_n = FeatureBuf_143;
         Mult_Buf[45].Weight_n = Wgt_9_143;
         Mult_Buf[46].Feature_n = FeatureBuf_144;
         Mult_Buf[46].Weight_n = Wgt_9_144;
         Mult_Buf[47].Feature_n = FeatureBuf_145;
         Mult_Buf[47].Weight_n = Wgt_9_145;
         Mult_Buf[48].Feature_n = FeatureBuf_146;
         Mult_Buf[48].Weight_n = Wgt_9_146;
         Mult_Buf[49].Feature_n = FeatureBuf_147;
         Mult_Buf[49].Weight_n = Wgt_9_147;
         Mult_Buf[50].Feature_n = FeatureBuf_148;
         Mult_Buf[50].Weight_n = Wgt_9_148;
         Mult_Buf[51].Feature_n = FeatureBuf_149;
         Mult_Buf[51].Weight_n = Wgt_9_149;
         Mult_Buf[52].Feature_n = FeatureBuf_150;
         Mult_Buf[52].Weight_n = Wgt_9_150;
         Mult_Buf[53].Feature_n = FeatureBuf_151;
         Mult_Buf[53].Weight_n = Wgt_9_151;
         Mult_Buf[54].Feature_n = FeatureBuf_152;
         Mult_Buf[54].Weight_n = Wgt_9_152;
         Mult_Buf[55].Feature_n = FeatureBuf_153;
         Mult_Buf[55].Weight_n = Wgt_9_153;
         Mult_Buf[56].Feature_n = FeatureBuf_154;
         Mult_Buf[56].Weight_n = Wgt_9_154;
         Mult_Buf[57].Feature_n = FeatureBuf_155;
         Mult_Buf[57].Weight_n = Wgt_9_155;
         Mult_Buf[58].Feature_n = FeatureBuf_156;
         Mult_Buf[58].Weight_n = Wgt_9_156;
         Mult_Buf[59].Feature_n = FeatureBuf_157;
         Mult_Buf[59].Weight_n = Wgt_9_157;
         Mult_Buf[60].Feature_n = FeatureBuf_158;
         Mult_Buf[60].Weight_n = Wgt_9_158;
         Mult_Buf[61].Feature_n = FeatureBuf_159;
         Mult_Buf[61].Weight_n = Wgt_9_159;
         Mult_Buf[62].Feature_n = FeatureBuf_160;
         Mult_Buf[62].Weight_n = Wgt_9_160;
         Mult_Buf[63].Feature_n = FeatureBuf_161;
         Mult_Buf[63].Weight_n = Wgt_9_161;
         Mult_Buf[64].Feature_n = FeatureBuf_162;
         Mult_Buf[64].Weight_n = Wgt_9_162;
         Mult_Buf[65].Feature_n = FeatureBuf_163;
         Mult_Buf[65].Weight_n = Wgt_9_163;
         Mult_Buf[66].Feature_n = FeatureBuf_164;
         Mult_Buf[66].Weight_n = Wgt_9_164;
         Mult_Buf[67].Feature_n = FeatureBuf_165;
         Mult_Buf[67].Weight_n = Wgt_9_165;
         Mult_Buf[68].Feature_n = FeatureBuf_166;
         Mult_Buf[68].Weight_n = Wgt_9_166;
         Mult_Buf[69].Feature_n = FeatureBuf_167;
         Mult_Buf[69].Weight_n = Wgt_9_167;
         Mult_Buf[70].Feature_n = FeatureBuf_168;
         Mult_Buf[70].Weight_n = Wgt_9_168;
         Mult_Buf[71].Feature_n = FeatureBuf_169;
         Mult_Buf[71].Weight_n = Wgt_9_169;
         Mult_Buf[72].Feature_n = FeatureBuf_170;
         Mult_Buf[72].Weight_n = Wgt_9_170;
         Mult_Buf[73].Feature_n = FeatureBuf_171;
         Mult_Buf[73].Weight_n = Wgt_9_171;
         Mult_Buf[74].Feature_n = FeatureBuf_172;
         Mult_Buf[74].Weight_n = Wgt_9_172;
         Mult_Buf[75].Feature_n = FeatureBuf_173;
         Mult_Buf[75].Weight_n = Wgt_9_173;
         Mult_Buf[76].Feature_n = FeatureBuf_174;
         Mult_Buf[76].Weight_n = Wgt_9_174;
         Mult_Buf[77].Feature_n = FeatureBuf_175;
         Mult_Buf[77].Weight_n = Wgt_9_175;
         Mult_Buf[78].Feature_n = FeatureBuf_176;
         Mult_Buf[78].Weight_n = Wgt_9_176;
         Mult_Buf[79].Feature_n = FeatureBuf_177;
         Mult_Buf[79].Weight_n = Wgt_9_177;
         Mult_Buf[80].Feature_n = FeatureBuf_178;
         Mult_Buf[80].Weight_n = Wgt_9_178;
         Mult_Buf[81].Feature_n = FeatureBuf_179;
         Mult_Buf[81].Weight_n = Wgt_9_179;
         Mult_Buf[82].Feature_n = FeatureBuf_180;
         Mult_Buf[82].Weight_n = Wgt_9_180;
         Mult_Buf[83].Feature_n = FeatureBuf_181;
         Mult_Buf[83].Weight_n = Wgt_9_181;
         Mult_Buf[84].Feature_n = FeatureBuf_182;
         Mult_Buf[84].Weight_n = Wgt_9_182;
         Mult_Buf[85].Feature_n = FeatureBuf_183;
         Mult_Buf[85].Weight_n = Wgt_9_183;
         Mult_Buf[86].Feature_n = FeatureBuf_184;
         Mult_Buf[86].Weight_n = Wgt_9_184;
         Mult_Buf[87].Feature_n = FeatureBuf_185;
         Mult_Buf[87].Weight_n = Wgt_9_185;
         Mult_Buf[88].Feature_n = FeatureBuf_186;
         Mult_Buf[88].Weight_n = Wgt_9_186;
         Mult_Buf[89].Feature_n = FeatureBuf_187;
         Mult_Buf[89].Weight_n = Wgt_9_187;
         Mult_Buf[90].Feature_n = FeatureBuf_188;
         Mult_Buf[90].Weight_n = Wgt_9_188;
         Mult_Buf[91].Feature_n = FeatureBuf_189;
         Mult_Buf[91].Weight_n = Wgt_9_189;
         Mult_Buf[92].Feature_n = FeatureBuf_190;
         Mult_Buf[92].Weight_n = Wgt_9_190;
         Mult_Buf[93].Feature_n = FeatureBuf_191;
         Mult_Buf[93].Weight_n = Wgt_9_191;
         Mult_Buf[94].Feature_n = FeatureBuf_192;
         Mult_Buf[94].Weight_n = Wgt_9_192;
         Mult_Buf[95].Feature_n = FeatureBuf_193;
         Mult_Buf[95].Weight_n = Wgt_9_193;
         Mult_Buf[96].Feature_n = FeatureBuf_194;
         Mult_Buf[96].Weight_n = Wgt_9_194;
         Mult_Buf[97].Feature_n = FeatureBuf_195;
         Mult_Buf[97].Weight_n = Wgt_9_195;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     //Collect Partial result form Adder
         Res_6_3_n = Part_Res;
     end
    76:begin
     nxt_state = 77;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_196;
         Mult_Buf[0].Weight_n = Wgt_9_196;
         Mult_Buf[1].Feature_n = FeatureBuf_197;
         Mult_Buf[1].Weight_n = Wgt_9_197;
         Mult_Buf[2].Feature_n = FeatureBuf_198;
         Mult_Buf[2].Weight_n = Wgt_9_198;
         Mult_Buf[3].Feature_n = FeatureBuf_199;
         Mult_Buf[3].Weight_n = Wgt_9_199;
         Mult_Buf[4].Feature_n = FeatureBuf_200;
         Mult_Buf[4].Weight_n = Wgt_9_200;
         Mult_Buf[5].Feature_n = FeatureBuf_201;
         Mult_Buf[5].Weight_n = Wgt_9_201;
         Mult_Buf[6].Feature_n = FeatureBuf_202;
         Mult_Buf[6].Weight_n = Wgt_9_202;
         Mult_Buf[7].Feature_n = FeatureBuf_203;
         Mult_Buf[7].Weight_n = Wgt_9_203;
         Mult_Buf[8].Feature_n = FeatureBuf_204;
         Mult_Buf[8].Weight_n = Wgt_9_204;
         Mult_Buf[9].Feature_n = FeatureBuf_205;
         Mult_Buf[9].Weight_n = Wgt_9_205;
         Mult_Buf[10].Feature_n = FeatureBuf_206;
         Mult_Buf[10].Weight_n = Wgt_9_206;
         Mult_Buf[11].Feature_n = FeatureBuf_207;
         Mult_Buf[11].Weight_n = Wgt_9_207;
         Mult_Buf[12].Feature_n = FeatureBuf_208;
         Mult_Buf[12].Weight_n = Wgt_9_208;
         Mult_Buf[13].Feature_n = FeatureBuf_209;
         Mult_Buf[13].Weight_n = Wgt_9_209;
         Mult_Buf[14].Feature_n = FeatureBuf_210;
         Mult_Buf[14].Weight_n = Wgt_9_210;
         Mult_Buf[15].Feature_n = FeatureBuf_211;
         Mult_Buf[15].Weight_n = Wgt_9_211;
         Mult_Buf[16].Feature_n = FeatureBuf_212;
         Mult_Buf[16].Weight_n = Wgt_9_212;
         Mult_Buf[17].Feature_n = FeatureBuf_213;
         Mult_Buf[17].Weight_n = Wgt_9_213;
         Mult_Buf[18].Feature_n = FeatureBuf_214;
         Mult_Buf[18].Weight_n = Wgt_9_214;
         Mult_Buf[19].Feature_n = FeatureBuf_215;
         Mult_Buf[19].Weight_n = Wgt_9_215;
         Mult_Buf[20].Feature_n = FeatureBuf_216;
         Mult_Buf[20].Weight_n = Wgt_9_216;
         Mult_Buf[21].Feature_n = FeatureBuf_217;
         Mult_Buf[21].Weight_n = Wgt_9_217;
         Mult_Buf[22].Feature_n = FeatureBuf_218;
         Mult_Buf[22].Weight_n = Wgt_9_218;
         Mult_Buf[23].Feature_n = FeatureBuf_219;
         Mult_Buf[23].Weight_n = Wgt_9_219;
         Mult_Buf[24].Feature_n = FeatureBuf_220;
         Mult_Buf[24].Weight_n = Wgt_9_220;
         Mult_Buf[25].Feature_n = FeatureBuf_221;
         Mult_Buf[25].Weight_n = Wgt_9_221;
         Mult_Buf[26].Feature_n = FeatureBuf_222;
         Mult_Buf[26].Weight_n = Wgt_9_222;
         Mult_Buf[27].Feature_n = FeatureBuf_223;
         Mult_Buf[27].Weight_n = Wgt_9_223;
         Mult_Buf[28].Feature_n = FeatureBuf_224;
         Mult_Buf[28].Weight_n = Wgt_9_224;
         Mult_Buf[29].Feature_n = FeatureBuf_225;
         Mult_Buf[29].Weight_n = Wgt_9_225;
         Mult_Buf[30].Feature_n = FeatureBuf_226;
         Mult_Buf[30].Weight_n = Wgt_9_226;
         Mult_Buf[31].Feature_n = FeatureBuf_227;
         Mult_Buf[31].Weight_n = Wgt_9_227;
         Mult_Buf[32].Feature_n = FeatureBuf_228;
         Mult_Buf[32].Weight_n = Wgt_9_228;
         Mult_Buf[33].Feature_n = FeatureBuf_229;
         Mult_Buf[33].Weight_n = Wgt_9_229;
         Mult_Buf[34].Feature_n = FeatureBuf_230;
         Mult_Buf[34].Weight_n = Wgt_9_230;
         Mult_Buf[35].Feature_n = FeatureBuf_231;
         Mult_Buf[35].Weight_n = Wgt_9_231;
         Mult_Buf[36].Feature_n = FeatureBuf_232;
         Mult_Buf[36].Weight_n = Wgt_9_232;
         Mult_Buf[37].Feature_n = FeatureBuf_233;
         Mult_Buf[37].Weight_n = Wgt_9_233;
         Mult_Buf[38].Feature_n = FeatureBuf_234;
         Mult_Buf[38].Weight_n = Wgt_9_234;
         Mult_Buf[39].Feature_n = FeatureBuf_235;
         Mult_Buf[39].Weight_n = Wgt_9_235;
         Mult_Buf[40].Feature_n = FeatureBuf_236;
         Mult_Buf[40].Weight_n = Wgt_9_236;
         Mult_Buf[41].Feature_n = FeatureBuf_237;
         Mult_Buf[41].Weight_n = Wgt_9_237;
         Mult_Buf[42].Feature_n = FeatureBuf_238;
         Mult_Buf[42].Weight_n = Wgt_9_238;
         Mult_Buf[43].Feature_n = FeatureBuf_239;
         Mult_Buf[43].Weight_n = Wgt_9_239;
         Mult_Buf[44].Feature_n = FeatureBuf_240;
         Mult_Buf[44].Weight_n = Wgt_9_240;
         Mult_Buf[45].Feature_n = FeatureBuf_241;
         Mult_Buf[45].Weight_n = Wgt_9_241;
         Mult_Buf[46].Feature_n = FeatureBuf_242;
         Mult_Buf[46].Weight_n = Wgt_9_242;
         Mult_Buf[47].Feature_n = FeatureBuf_243;
         Mult_Buf[47].Weight_n = Wgt_9_243;
         Mult_Buf[48].Feature_n = FeatureBuf_244;
         Mult_Buf[48].Weight_n = Wgt_9_244;
         Mult_Buf[49].Feature_n = FeatureBuf_245;
         Mult_Buf[49].Weight_n = Wgt_9_245;
         Mult_Buf[50].Feature_n = FeatureBuf_246;
         Mult_Buf[50].Weight_n = Wgt_9_246;
         Mult_Buf[51].Feature_n = FeatureBuf_247;
         Mult_Buf[51].Weight_n = Wgt_9_247;
         Mult_Buf[52].Feature_n = FeatureBuf_248;
         Mult_Buf[52].Weight_n = Wgt_9_248;
         Mult_Buf[53].Feature_n = FeatureBuf_249;
         Mult_Buf[53].Weight_n = Wgt_9_249;
         Mult_Buf[54].Feature_n = FeatureBuf_250;
         Mult_Buf[54].Weight_n = Wgt_9_250;
         Mult_Buf[55].Feature_n = FeatureBuf_251;
         Mult_Buf[55].Weight_n = Wgt_9_251;
         Mult_Buf[56].Feature_n = FeatureBuf_252;
         Mult_Buf[56].Weight_n = Wgt_9_252;
         Mult_Buf[57].Feature_n = FeatureBuf_253;
         Mult_Buf[57].Weight_n = Wgt_9_253;
         Mult_Buf[58].Feature_n = FeatureBuf_254;
         Mult_Buf[58].Weight_n = Wgt_9_254;
         Mult_Buf[59].Feature_n = FeatureBuf_255;
         Mult_Buf[59].Weight_n = Wgt_9_255;
         Mult_Buf[60].Feature_n = FeatureBuf_256;
         Mult_Buf[60].Weight_n = Wgt_9_256;
         Mult_Buf[61].Feature_n = FeatureBuf_257;
         Mult_Buf[61].Weight_n = Wgt_9_257;
         Mult_Buf[62].Feature_n = FeatureBuf_258;
         Mult_Buf[62].Weight_n = Wgt_9_258;
         Mult_Buf[63].Feature_n = FeatureBuf_259;
         Mult_Buf[63].Weight_n = Wgt_9_259;
         Mult_Buf[64].Feature_n = FeatureBuf_260;
         Mult_Buf[64].Weight_n = Wgt_9_260;
         Mult_Buf[65].Feature_n = FeatureBuf_261;
         Mult_Buf[65].Weight_n = Wgt_9_261;
         Mult_Buf[66].Feature_n = FeatureBuf_262;
         Mult_Buf[66].Weight_n = Wgt_9_262;
         Mult_Buf[67].Feature_n = FeatureBuf_263;
         Mult_Buf[67].Weight_n = Wgt_9_263;
         Mult_Buf[68].Feature_n = FeatureBuf_264;
         Mult_Buf[68].Weight_n = Wgt_9_264;
         Mult_Buf[69].Feature_n = FeatureBuf_265;
         Mult_Buf[69].Weight_n = Wgt_9_265;
         Mult_Buf[70].Feature_n = FeatureBuf_266;
         Mult_Buf[70].Weight_n = Wgt_9_266;
         Mult_Buf[71].Feature_n = FeatureBuf_267;
         Mult_Buf[71].Weight_n = Wgt_9_267;
         Mult_Buf[72].Feature_n = FeatureBuf_268;
         Mult_Buf[72].Weight_n = Wgt_9_268;
         Mult_Buf[73].Feature_n = FeatureBuf_269;
         Mult_Buf[73].Weight_n = Wgt_9_269;
         Mult_Buf[74].Feature_n = FeatureBuf_270;
         Mult_Buf[74].Weight_n = Wgt_9_270;
         Mult_Buf[75].Feature_n = FeatureBuf_271;
         Mult_Buf[75].Weight_n = Wgt_9_271;
         Mult_Buf[76].Feature_n = FeatureBuf_272;
         Mult_Buf[76].Weight_n = Wgt_9_272;
         Mult_Buf[77].Feature_n = FeatureBuf_273;
         Mult_Buf[77].Weight_n = Wgt_9_273;
         Mult_Buf[78].Feature_n = FeatureBuf_274;
         Mult_Buf[78].Weight_n = Wgt_9_274;
         Mult_Buf[79].Feature_n = FeatureBuf_275;
         Mult_Buf[79].Weight_n = Wgt_9_275;
         Mult_Buf[80].Feature_n = FeatureBuf_276;
         Mult_Buf[80].Weight_n = Wgt_9_276;
         Mult_Buf[81].Feature_n = FeatureBuf_277;
         Mult_Buf[81].Weight_n = Wgt_9_277;
         Mult_Buf[82].Feature_n = FeatureBuf_278;
         Mult_Buf[82].Weight_n = Wgt_9_278;
         Mult_Buf[83].Feature_n = FeatureBuf_279;
         Mult_Buf[83].Weight_n = Wgt_9_279;
         Mult_Buf[84].Feature_n = FeatureBuf_280;
         Mult_Buf[84].Weight_n = Wgt_9_280;
         Mult_Buf[85].Feature_n = FeatureBuf_281;
         Mult_Buf[85].Weight_n = Wgt_9_281;
         Mult_Buf[86].Feature_n = FeatureBuf_282;
         Mult_Buf[86].Weight_n = Wgt_9_282;
         Mult_Buf[87].Feature_n = FeatureBuf_283;
         Mult_Buf[87].Weight_n = Wgt_9_283;
         Mult_Buf[88].Feature_n = FeatureBuf_284;
         Mult_Buf[88].Weight_n = Wgt_9_284;
         Mult_Buf[89].Feature_n = FeatureBuf_285;
         Mult_Buf[89].Weight_n = Wgt_9_285;
         Mult_Buf[90].Feature_n = FeatureBuf_286;
         Mult_Buf[90].Weight_n = Wgt_9_286;
         Mult_Buf[91].Feature_n = FeatureBuf_287;
         Mult_Buf[91].Weight_n = Wgt_9_287;
         Mult_Buf[92].Feature_n = FeatureBuf_288;
         Mult_Buf[92].Weight_n = Wgt_9_288;
         Mult_Buf[93].Feature_n = FeatureBuf_289;
         Mult_Buf[93].Weight_n = Wgt_9_289;
         Mult_Buf[94].Feature_n = FeatureBuf_290;
         Mult_Buf[94].Weight_n = Wgt_9_290;
         Mult_Buf[95].Feature_n = FeatureBuf_291;
         Mult_Buf[95].Weight_n = Wgt_9_291;
         Mult_Buf[96].Feature_n = FeatureBuf_292;
         Mult_Buf[96].Weight_n = Wgt_9_292;
         Mult_Buf[97].Feature_n = FeatureBuf_293;
         Mult_Buf[97].Weight_n = Wgt_9_293;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     //Collect Partial result form Adder
         Res_6_4_n = Part_Res;
     end
    77:begin
     nxt_state = 78;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_294;
         Mult_Buf[0].Weight_n = Wgt_9_294;
         Mult_Buf[1].Feature_n = FeatureBuf_295;
         Mult_Buf[1].Weight_n = Wgt_9_295;
         Mult_Buf[2].Feature_n = FeatureBuf_296;
         Mult_Buf[2].Weight_n = Wgt_9_296;
         Mult_Buf[3].Feature_n = FeatureBuf_297;
         Mult_Buf[3].Weight_n = Wgt_9_297;
         Mult_Buf[4].Feature_n = FeatureBuf_298;
         Mult_Buf[4].Weight_n = Wgt_9_298;
         Mult_Buf[5].Feature_n = FeatureBuf_299;
         Mult_Buf[5].Weight_n = Wgt_9_299;
         Mult_Buf[6].Feature_n = FeatureBuf_300;
         Mult_Buf[6].Weight_n = Wgt_9_300;
         Mult_Buf[7].Feature_n = FeatureBuf_301;
         Mult_Buf[7].Weight_n = Wgt_9_301;
         Mult_Buf[8].Feature_n = FeatureBuf_302;
         Mult_Buf[8].Weight_n = Wgt_9_302;
         Mult_Buf[9].Feature_n = FeatureBuf_303;
         Mult_Buf[9].Weight_n = Wgt_9_303;
         Mult_Buf[10].Feature_n = FeatureBuf_304;
         Mult_Buf[10].Weight_n = Wgt_9_304;
         Mult_Buf[11].Feature_n = FeatureBuf_305;
         Mult_Buf[11].Weight_n = Wgt_9_305;
         Mult_Buf[12].Feature_n = FeatureBuf_306;
         Mult_Buf[12].Weight_n = Wgt_9_306;
         Mult_Buf[13].Feature_n = FeatureBuf_307;
         Mult_Buf[13].Weight_n = Wgt_9_307;
         Mult_Buf[14].Feature_n = FeatureBuf_308;
         Mult_Buf[14].Weight_n = Wgt_9_308;
         Mult_Buf[15].Feature_n = FeatureBuf_309;
         Mult_Buf[15].Weight_n = Wgt_9_309;
         Mult_Buf[16].Feature_n = FeatureBuf_310;
         Mult_Buf[16].Weight_n = Wgt_9_310;
         Mult_Buf[17].Feature_n = FeatureBuf_311;
         Mult_Buf[17].Weight_n = Wgt_9_311;
         Mult_Buf[18].Feature_n = FeatureBuf_312;
         Mult_Buf[18].Weight_n = Wgt_9_312;
         Mult_Buf[19].Feature_n = FeatureBuf_313;
         Mult_Buf[19].Weight_n = Wgt_9_313;
         Mult_Buf[20].Feature_n = FeatureBuf_314;
         Mult_Buf[20].Weight_n = Wgt_9_314;
         Mult_Buf[21].Feature_n = FeatureBuf_315;
         Mult_Buf[21].Weight_n = Wgt_9_315;
         Mult_Buf[22].Feature_n = FeatureBuf_316;
         Mult_Buf[22].Weight_n = Wgt_9_316;
         Mult_Buf[23].Feature_n = FeatureBuf_317;
         Mult_Buf[23].Weight_n = Wgt_9_317;
         Mult_Buf[24].Feature_n = FeatureBuf_318;
         Mult_Buf[24].Weight_n = Wgt_9_318;
         Mult_Buf[25].Feature_n = FeatureBuf_319;
         Mult_Buf[25].Weight_n = Wgt_9_319;
         Mult_Buf[26].Feature_n = FeatureBuf_320;
         Mult_Buf[26].Weight_n = Wgt_9_320;
         Mult_Buf[27].Feature_n = FeatureBuf_321;
         Mult_Buf[27].Weight_n = Wgt_9_321;
         Mult_Buf[28].Feature_n = FeatureBuf_322;
         Mult_Buf[28].Weight_n = Wgt_9_322;
         Mult_Buf[29].Feature_n = FeatureBuf_323;
         Mult_Buf[29].Weight_n = Wgt_9_323;
         Mult_Buf[30].Feature_n = FeatureBuf_324;
         Mult_Buf[30].Weight_n = Wgt_9_324;
         Mult_Buf[31].Feature_n = FeatureBuf_325;
         Mult_Buf[31].Weight_n = Wgt_9_325;
         Mult_Buf[32].Feature_n = FeatureBuf_326;
         Mult_Buf[32].Weight_n = Wgt_9_326;
         Mult_Buf[33].Feature_n = FeatureBuf_327;
         Mult_Buf[33].Weight_n = Wgt_9_327;
         Mult_Buf[34].Feature_n = FeatureBuf_328;
         Mult_Buf[34].Weight_n = Wgt_9_328;
         Mult_Buf[35].Feature_n = FeatureBuf_329;
         Mult_Buf[35].Weight_n = Wgt_9_329;
         Mult_Buf[36].Feature_n = FeatureBuf_330;
         Mult_Buf[36].Weight_n = Wgt_9_330;
         Mult_Buf[37].Feature_n = FeatureBuf_331;
         Mult_Buf[37].Weight_n = Wgt_9_331;
         Mult_Buf[38].Feature_n = FeatureBuf_332;
         Mult_Buf[38].Weight_n = Wgt_9_332;
         Mult_Buf[39].Feature_n = FeatureBuf_333;
         Mult_Buf[39].Weight_n = Wgt_9_333;
         Mult_Buf[40].Feature_n = FeatureBuf_334;
         Mult_Buf[40].Weight_n = Wgt_9_334;
         Mult_Buf[41].Feature_n = FeatureBuf_335;
         Mult_Buf[41].Weight_n = Wgt_9_335;
         Mult_Buf[42].Feature_n = FeatureBuf_336;
         Mult_Buf[42].Weight_n = Wgt_9_336;
         Mult_Buf[43].Feature_n = FeatureBuf_337;
         Mult_Buf[43].Weight_n = Wgt_9_337;
         Mult_Buf[44].Feature_n = FeatureBuf_338;
         Mult_Buf[44].Weight_n = Wgt_9_338;
         Mult_Buf[45].Feature_n = FeatureBuf_339;
         Mult_Buf[45].Weight_n = Wgt_9_339;
         Mult_Buf[46].Feature_n = FeatureBuf_340;
         Mult_Buf[46].Weight_n = Wgt_9_340;
         Mult_Buf[47].Feature_n = FeatureBuf_341;
         Mult_Buf[47].Weight_n = Wgt_9_341;
         Mult_Buf[48].Feature_n = FeatureBuf_342;
         Mult_Buf[48].Weight_n = Wgt_9_342;
         Mult_Buf[49].Feature_n = FeatureBuf_343;
         Mult_Buf[49].Weight_n = Wgt_9_343;
         Mult_Buf[50].Feature_n = FeatureBuf_344;
         Mult_Buf[50].Weight_n = Wgt_9_344;
         Mult_Buf[51].Feature_n = FeatureBuf_345;
         Mult_Buf[51].Weight_n = Wgt_9_345;
         Mult_Buf[52].Feature_n = FeatureBuf_346;
         Mult_Buf[52].Weight_n = Wgt_9_346;
         Mult_Buf[53].Feature_n = FeatureBuf_347;
         Mult_Buf[53].Weight_n = Wgt_9_347;
         Mult_Buf[54].Feature_n = FeatureBuf_348;
         Mult_Buf[54].Weight_n = Wgt_9_348;
         Mult_Buf[55].Feature_n = FeatureBuf_349;
         Mult_Buf[55].Weight_n = Wgt_9_349;
         Mult_Buf[56].Feature_n = FeatureBuf_350;
         Mult_Buf[56].Weight_n = Wgt_9_350;
         Mult_Buf[57].Feature_n = FeatureBuf_351;
         Mult_Buf[57].Weight_n = Wgt_9_351;
         Mult_Buf[58].Feature_n = FeatureBuf_352;
         Mult_Buf[58].Weight_n = Wgt_9_352;
         Mult_Buf[59].Feature_n = FeatureBuf_353;
         Mult_Buf[59].Weight_n = Wgt_9_353;
         Mult_Buf[60].Feature_n = FeatureBuf_354;
         Mult_Buf[60].Weight_n = Wgt_9_354;
         Mult_Buf[61].Feature_n = FeatureBuf_355;
         Mult_Buf[61].Weight_n = Wgt_9_355;
         Mult_Buf[62].Feature_n = FeatureBuf_356;
         Mult_Buf[62].Weight_n = Wgt_9_356;
         Mult_Buf[63].Feature_n = FeatureBuf_357;
         Mult_Buf[63].Weight_n = Wgt_9_357;
         Mult_Buf[64].Feature_n = FeatureBuf_358;
         Mult_Buf[64].Weight_n = Wgt_9_358;
         Mult_Buf[65].Feature_n = FeatureBuf_359;
         Mult_Buf[65].Weight_n = Wgt_9_359;
         Mult_Buf[66].Feature_n = FeatureBuf_360;
         Mult_Buf[66].Weight_n = Wgt_9_360;
         Mult_Buf[67].Feature_n = FeatureBuf_361;
         Mult_Buf[67].Weight_n = Wgt_9_361;
         Mult_Buf[68].Feature_n = FeatureBuf_362;
         Mult_Buf[68].Weight_n = Wgt_9_362;
         Mult_Buf[69].Feature_n = FeatureBuf_363;
         Mult_Buf[69].Weight_n = Wgt_9_363;
         Mult_Buf[70].Feature_n = FeatureBuf_364;
         Mult_Buf[70].Weight_n = Wgt_9_364;
         Mult_Buf[71].Feature_n = FeatureBuf_365;
         Mult_Buf[71].Weight_n = Wgt_9_365;
         Mult_Buf[72].Feature_n = FeatureBuf_366;
         Mult_Buf[72].Weight_n = Wgt_9_366;
         Mult_Buf[73].Feature_n = FeatureBuf_367;
         Mult_Buf[73].Weight_n = Wgt_9_367;
         Mult_Buf[74].Feature_n = FeatureBuf_368;
         Mult_Buf[74].Weight_n = Wgt_9_368;
         Mult_Buf[75].Feature_n = FeatureBuf_369;
         Mult_Buf[75].Weight_n = Wgt_9_369;
         Mult_Buf[76].Feature_n = FeatureBuf_370;
         Mult_Buf[76].Weight_n = Wgt_9_370;
         Mult_Buf[77].Feature_n = FeatureBuf_371;
         Mult_Buf[77].Weight_n = Wgt_9_371;
         Mult_Buf[78].Feature_n = FeatureBuf_372;
         Mult_Buf[78].Weight_n = Wgt_9_372;
         Mult_Buf[79].Feature_n = FeatureBuf_373;
         Mult_Buf[79].Weight_n = Wgt_9_373;
         Mult_Buf[80].Feature_n = FeatureBuf_374;
         Mult_Buf[80].Weight_n = Wgt_9_374;
         Mult_Buf[81].Feature_n = FeatureBuf_375;
         Mult_Buf[81].Weight_n = Wgt_9_375;
         Mult_Buf[82].Feature_n = FeatureBuf_376;
         Mult_Buf[82].Weight_n = Wgt_9_376;
         Mult_Buf[83].Feature_n = FeatureBuf_377;
         Mult_Buf[83].Weight_n = Wgt_9_377;
         Mult_Buf[84].Feature_n = FeatureBuf_378;
         Mult_Buf[84].Weight_n = Wgt_9_378;
         Mult_Buf[85].Feature_n = FeatureBuf_379;
         Mult_Buf[85].Weight_n = Wgt_9_379;
         Mult_Buf[86].Feature_n = FeatureBuf_380;
         Mult_Buf[86].Weight_n = Wgt_9_380;
         Mult_Buf[87].Feature_n = FeatureBuf_381;
         Mult_Buf[87].Weight_n = Wgt_9_381;
         Mult_Buf[88].Feature_n = FeatureBuf_382;
         Mult_Buf[88].Weight_n = Wgt_9_382;
         Mult_Buf[89].Feature_n = FeatureBuf_383;
         Mult_Buf[89].Weight_n = Wgt_9_383;
         Mult_Buf[90].Feature_n = FeatureBuf_384;
         Mult_Buf[90].Weight_n = Wgt_9_384;
         Mult_Buf[91].Feature_n = FeatureBuf_385;
         Mult_Buf[91].Weight_n = Wgt_9_385;
         Mult_Buf[92].Feature_n = FeatureBuf_386;
         Mult_Buf[92].Weight_n = Wgt_9_386;
         Mult_Buf[93].Feature_n = FeatureBuf_387;
         Mult_Buf[93].Weight_n = Wgt_9_387;
         Mult_Buf[94].Feature_n = FeatureBuf_388;
         Mult_Buf[94].Weight_n = Wgt_9_388;
         Mult_Buf[95].Feature_n = FeatureBuf_389;
         Mult_Buf[95].Weight_n = Wgt_9_389;
         Mult_Buf[96].Feature_n = FeatureBuf_390;
         Mult_Buf[96].Weight_n = Wgt_9_390;
         Mult_Buf[97].Feature_n = FeatureBuf_391;
         Mult_Buf[97].Weight_n = Wgt_9_391;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     //Collect Partial result form Adder
         Res_6_5_n = Part_Res;
     //Collect result from final Adder
         Res5_n = Final_Res;
     end
    78:begin
     nxt_state = 79;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_392;
         Mult_Buf[0].Weight_n = Wgt_9_392;
         Mult_Buf[1].Feature_n = FeatureBuf_393;
         Mult_Buf[1].Weight_n = Wgt_9_393;
         Mult_Buf[2].Feature_n = FeatureBuf_394;
         Mult_Buf[2].Weight_n = Wgt_9_394;
         Mult_Buf[3].Feature_n = FeatureBuf_395;
         Mult_Buf[3].Weight_n = Wgt_9_395;
         Mult_Buf[4].Feature_n = FeatureBuf_396;
         Mult_Buf[4].Weight_n = Wgt_9_396;
         Mult_Buf[5].Feature_n = FeatureBuf_397;
         Mult_Buf[5].Weight_n = Wgt_9_397;
         Mult_Buf[6].Feature_n = FeatureBuf_398;
         Mult_Buf[6].Weight_n = Wgt_9_398;
         Mult_Buf[7].Feature_n = FeatureBuf_399;
         Mult_Buf[7].Weight_n = Wgt_9_399;
         Mult_Buf[8].Feature_n = FeatureBuf_400;
         Mult_Buf[8].Weight_n = Wgt_9_400;
         Mult_Buf[9].Feature_n = FeatureBuf_401;
         Mult_Buf[9].Weight_n = Wgt_9_401;
         Mult_Buf[10].Feature_n = FeatureBuf_402;
         Mult_Buf[10].Weight_n = Wgt_9_402;
         Mult_Buf[11].Feature_n = FeatureBuf_403;
         Mult_Buf[11].Weight_n = Wgt_9_403;
         Mult_Buf[12].Feature_n = FeatureBuf_404;
         Mult_Buf[12].Weight_n = Wgt_9_404;
         Mult_Buf[13].Feature_n = FeatureBuf_405;
         Mult_Buf[13].Weight_n = Wgt_9_405;
         Mult_Buf[14].Feature_n = FeatureBuf_406;
         Mult_Buf[14].Weight_n = Wgt_9_406;
         Mult_Buf[15].Feature_n = FeatureBuf_407;
         Mult_Buf[15].Weight_n = Wgt_9_407;
         Mult_Buf[16].Feature_n = FeatureBuf_408;
         Mult_Buf[16].Weight_n = Wgt_9_408;
         Mult_Buf[17].Feature_n = FeatureBuf_409;
         Mult_Buf[17].Weight_n = Wgt_9_409;
         Mult_Buf[18].Feature_n = FeatureBuf_410;
         Mult_Buf[18].Weight_n = Wgt_9_410;
         Mult_Buf[19].Feature_n = FeatureBuf_411;
         Mult_Buf[19].Weight_n = Wgt_9_411;
         Mult_Buf[20].Feature_n = FeatureBuf_412;
         Mult_Buf[20].Weight_n = Wgt_9_412;
         Mult_Buf[21].Feature_n = FeatureBuf_413;
         Mult_Buf[21].Weight_n = Wgt_9_413;
         Mult_Buf[22].Feature_n = FeatureBuf_414;
         Mult_Buf[22].Weight_n = Wgt_9_414;
         Mult_Buf[23].Feature_n = FeatureBuf_415;
         Mult_Buf[23].Weight_n = Wgt_9_415;
         Mult_Buf[24].Feature_n = FeatureBuf_416;
         Mult_Buf[24].Weight_n = Wgt_9_416;
         Mult_Buf[25].Feature_n = FeatureBuf_417;
         Mult_Buf[25].Weight_n = Wgt_9_417;
         Mult_Buf[26].Feature_n = FeatureBuf_418;
         Mult_Buf[26].Weight_n = Wgt_9_418;
         Mult_Buf[27].Feature_n = FeatureBuf_419;
         Mult_Buf[27].Weight_n = Wgt_9_419;
         Mult_Buf[28].Feature_n = FeatureBuf_420;
         Mult_Buf[28].Weight_n = Wgt_9_420;
         Mult_Buf[29].Feature_n = FeatureBuf_421;
         Mult_Buf[29].Weight_n = Wgt_9_421;
         Mult_Buf[30].Feature_n = FeatureBuf_422;
         Mult_Buf[30].Weight_n = Wgt_9_422;
         Mult_Buf[31].Feature_n = FeatureBuf_423;
         Mult_Buf[31].Weight_n = Wgt_9_423;
         Mult_Buf[32].Feature_n = FeatureBuf_424;
         Mult_Buf[32].Weight_n = Wgt_9_424;
         Mult_Buf[33].Feature_n = FeatureBuf_425;
         Mult_Buf[33].Weight_n = Wgt_9_425;
         Mult_Buf[34].Feature_n = FeatureBuf_426;
         Mult_Buf[34].Weight_n = Wgt_9_426;
         Mult_Buf[35].Feature_n = FeatureBuf_427;
         Mult_Buf[35].Weight_n = Wgt_9_427;
         Mult_Buf[36].Feature_n = FeatureBuf_428;
         Mult_Buf[36].Weight_n = Wgt_9_428;
         Mult_Buf[37].Feature_n = FeatureBuf_429;
         Mult_Buf[37].Weight_n = Wgt_9_429;
         Mult_Buf[38].Feature_n = FeatureBuf_430;
         Mult_Buf[38].Weight_n = Wgt_9_430;
         Mult_Buf[39].Feature_n = FeatureBuf_431;
         Mult_Buf[39].Weight_n = Wgt_9_431;
         Mult_Buf[40].Feature_n = FeatureBuf_432;
         Mult_Buf[40].Weight_n = Wgt_9_432;
         Mult_Buf[41].Feature_n = FeatureBuf_433;
         Mult_Buf[41].Weight_n = Wgt_9_433;
         Mult_Buf[42].Feature_n = FeatureBuf_434;
         Mult_Buf[42].Weight_n = Wgt_9_434;
         Mult_Buf[43].Feature_n = FeatureBuf_435;
         Mult_Buf[43].Weight_n = Wgt_9_435;
         Mult_Buf[44].Feature_n = FeatureBuf_436;
         Mult_Buf[44].Weight_n = Wgt_9_436;
         Mult_Buf[45].Feature_n = FeatureBuf_437;
         Mult_Buf[45].Weight_n = Wgt_9_437;
         Mult_Buf[46].Feature_n = FeatureBuf_438;
         Mult_Buf[46].Weight_n = Wgt_9_438;
         Mult_Buf[47].Feature_n = FeatureBuf_439;
         Mult_Buf[47].Weight_n = Wgt_9_439;
         Mult_Buf[48].Feature_n = FeatureBuf_440;
         Mult_Buf[48].Weight_n = Wgt_9_440;
         Mult_Buf[49].Feature_n = FeatureBuf_441;
         Mult_Buf[49].Weight_n = Wgt_9_441;
         Mult_Buf[50].Feature_n = FeatureBuf_442;
         Mult_Buf[50].Weight_n = Wgt_9_442;
         Mult_Buf[51].Feature_n = FeatureBuf_443;
         Mult_Buf[51].Weight_n = Wgt_9_443;
         Mult_Buf[52].Feature_n = FeatureBuf_444;
         Mult_Buf[52].Weight_n = Wgt_9_444;
         Mult_Buf[53].Feature_n = FeatureBuf_445;
         Mult_Buf[53].Weight_n = Wgt_9_445;
         Mult_Buf[54].Feature_n = FeatureBuf_446;
         Mult_Buf[54].Weight_n = Wgt_9_446;
         Mult_Buf[55].Feature_n = FeatureBuf_447;
         Mult_Buf[55].Weight_n = Wgt_9_447;
         Mult_Buf[56].Feature_n = FeatureBuf_448;
         Mult_Buf[56].Weight_n = Wgt_9_448;
         Mult_Buf[57].Feature_n = FeatureBuf_449;
         Mult_Buf[57].Weight_n = Wgt_9_449;
         Mult_Buf[58].Feature_n = FeatureBuf_450;
         Mult_Buf[58].Weight_n = Wgt_9_450;
         Mult_Buf[59].Feature_n = FeatureBuf_451;
         Mult_Buf[59].Weight_n = Wgt_9_451;
         Mult_Buf[60].Feature_n = FeatureBuf_452;
         Mult_Buf[60].Weight_n = Wgt_9_452;
         Mult_Buf[61].Feature_n = FeatureBuf_453;
         Mult_Buf[61].Weight_n = Wgt_9_453;
         Mult_Buf[62].Feature_n = FeatureBuf_454;
         Mult_Buf[62].Weight_n = Wgt_9_454;
         Mult_Buf[63].Feature_n = FeatureBuf_455;
         Mult_Buf[63].Weight_n = Wgt_9_455;
         Mult_Buf[64].Feature_n = FeatureBuf_456;
         Mult_Buf[64].Weight_n = Wgt_9_456;
         Mult_Buf[65].Feature_n = FeatureBuf_457;
         Mult_Buf[65].Weight_n = Wgt_9_457;
         Mult_Buf[66].Feature_n = FeatureBuf_458;
         Mult_Buf[66].Weight_n = Wgt_9_458;
         Mult_Buf[67].Feature_n = FeatureBuf_459;
         Mult_Buf[67].Weight_n = Wgt_9_459;
         Mult_Buf[68].Feature_n = FeatureBuf_460;
         Mult_Buf[68].Weight_n = Wgt_9_460;
         Mult_Buf[69].Feature_n = FeatureBuf_461;
         Mult_Buf[69].Weight_n = Wgt_9_461;
         Mult_Buf[70].Feature_n = FeatureBuf_462;
         Mult_Buf[70].Weight_n = Wgt_9_462;
         Mult_Buf[71].Feature_n = FeatureBuf_463;
         Mult_Buf[71].Weight_n = Wgt_9_463;
         Mult_Buf[72].Feature_n = FeatureBuf_464;
         Mult_Buf[72].Weight_n = Wgt_9_464;
         Mult_Buf[73].Feature_n = FeatureBuf_465;
         Mult_Buf[73].Weight_n = Wgt_9_465;
         Mult_Buf[74].Feature_n = FeatureBuf_466;
         Mult_Buf[74].Weight_n = Wgt_9_466;
         Mult_Buf[75].Feature_n = FeatureBuf_467;
         Mult_Buf[75].Weight_n = Wgt_9_467;
         Mult_Buf[76].Feature_n = FeatureBuf_468;
         Mult_Buf[76].Weight_n = Wgt_9_468;
         Mult_Buf[77].Feature_n = FeatureBuf_469;
         Mult_Buf[77].Weight_n = Wgt_9_469;
         Mult_Buf[78].Feature_n = FeatureBuf_470;
         Mult_Buf[78].Weight_n = Wgt_9_470;
         Mult_Buf[79].Feature_n = FeatureBuf_471;
         Mult_Buf[79].Weight_n = Wgt_9_471;
         Mult_Buf[80].Feature_n = FeatureBuf_472;
         Mult_Buf[80].Weight_n = Wgt_9_472;
         Mult_Buf[81].Feature_n = FeatureBuf_473;
         Mult_Buf[81].Weight_n = Wgt_9_473;
         Mult_Buf[82].Feature_n = FeatureBuf_474;
         Mult_Buf[82].Weight_n = Wgt_9_474;
         Mult_Buf[83].Feature_n = FeatureBuf_475;
         Mult_Buf[83].Weight_n = Wgt_9_475;
         Mult_Buf[84].Feature_n = FeatureBuf_476;
         Mult_Buf[84].Weight_n = Wgt_9_476;
         Mult_Buf[85].Feature_n = FeatureBuf_477;
         Mult_Buf[85].Weight_n = Wgt_9_477;
         Mult_Buf[86].Feature_n = FeatureBuf_478;
         Mult_Buf[86].Weight_n = Wgt_9_478;
         Mult_Buf[87].Feature_n = FeatureBuf_479;
         Mult_Buf[87].Weight_n = Wgt_9_479;
         Mult_Buf[88].Feature_n = FeatureBuf_480;
         Mult_Buf[88].Weight_n = Wgt_9_480;
         Mult_Buf[89].Feature_n = FeatureBuf_481;
         Mult_Buf[89].Weight_n = Wgt_9_481;
         Mult_Buf[90].Feature_n = FeatureBuf_482;
         Mult_Buf[90].Weight_n = Wgt_9_482;
         Mult_Buf[91].Feature_n = FeatureBuf_483;
         Mult_Buf[91].Weight_n = Wgt_9_483;
         Mult_Buf[92].Feature_n = FeatureBuf_484;
         Mult_Buf[92].Weight_n = Wgt_9_484;
         Mult_Buf[93].Feature_n = FeatureBuf_485;
         Mult_Buf[93].Weight_n = Wgt_9_485;
         Mult_Buf[94].Feature_n = FeatureBuf_486;
         Mult_Buf[94].Weight_n = Wgt_9_486;
         Mult_Buf[95].Feature_n = FeatureBuf_487;
         Mult_Buf[95].Weight_n = Wgt_9_487;
         Mult_Buf[96].Feature_n = FeatureBuf_488;
         Mult_Buf[96].Weight_n = Wgt_9_488;
         Mult_Buf[97].Feature_n = FeatureBuf_489;
         Mult_Buf[97].Weight_n = Wgt_9_489;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     //Collect Partial result form Adder
         Res_6_6_n = Part_Res;
     end
    79:begin
     nxt_state = 80;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_490;
         Mult_Buf[0].Weight_n = Wgt_9_490;
         Mult_Buf[1].Feature_n = FeatureBuf_491;
         Mult_Buf[1].Weight_n = Wgt_9_491;
         Mult_Buf[2].Feature_n = FeatureBuf_492;
         Mult_Buf[2].Weight_n = Wgt_9_492;
         Mult_Buf[3].Feature_n = FeatureBuf_493;
         Mult_Buf[3].Weight_n = Wgt_9_493;
         Mult_Buf[4].Feature_n = FeatureBuf_494;
         Mult_Buf[4].Weight_n = Wgt_9_494;
         Mult_Buf[5].Feature_n = FeatureBuf_495;
         Mult_Buf[5].Weight_n = Wgt_9_495;
         Mult_Buf[6].Feature_n = FeatureBuf_496;
         Mult_Buf[6].Weight_n = Wgt_9_496;
         Mult_Buf[7].Feature_n = FeatureBuf_497;
         Mult_Buf[7].Weight_n = Wgt_9_497;
         Mult_Buf[8].Feature_n = FeatureBuf_498;
         Mult_Buf[8].Weight_n = Wgt_9_498;
         Mult_Buf[9].Feature_n = FeatureBuf_499;
         Mult_Buf[9].Weight_n = Wgt_9_499;
         Mult_Buf[10].Feature_n = FeatureBuf_500;
         Mult_Buf[10].Weight_n = Wgt_9_500;
         Mult_Buf[11].Feature_n = FeatureBuf_501;
         Mult_Buf[11].Weight_n = Wgt_9_501;
         Mult_Buf[12].Feature_n = FeatureBuf_502;
         Mult_Buf[12].Weight_n = Wgt_9_502;
         Mult_Buf[13].Feature_n = FeatureBuf_503;
         Mult_Buf[13].Weight_n = Wgt_9_503;
         Mult_Buf[14].Feature_n = FeatureBuf_504;
         Mult_Buf[14].Weight_n = Wgt_9_504;
         Mult_Buf[15].Feature_n = FeatureBuf_505;
         Mult_Buf[15].Weight_n = Wgt_9_505;
         Mult_Buf[16].Feature_n = FeatureBuf_506;
         Mult_Buf[16].Weight_n = Wgt_9_506;
         Mult_Buf[17].Feature_n = FeatureBuf_507;
         Mult_Buf[17].Weight_n = Wgt_9_507;
         Mult_Buf[18].Feature_n = FeatureBuf_508;
         Mult_Buf[18].Weight_n = Wgt_9_508;
         Mult_Buf[19].Feature_n = FeatureBuf_509;
         Mult_Buf[19].Weight_n = Wgt_9_509;
         Mult_Buf[20].Feature_n = FeatureBuf_510;
         Mult_Buf[20].Weight_n = Wgt_9_510;
         Mult_Buf[21].Feature_n = FeatureBuf_511;
         Mult_Buf[21].Weight_n = Wgt_9_511;
         Mult_Buf[22].Feature_n = FeatureBuf_512;
         Mult_Buf[22].Weight_n = Wgt_9_512;
         Mult_Buf[23].Feature_n = FeatureBuf_513;
         Mult_Buf[23].Weight_n = Wgt_9_513;
         Mult_Buf[24].Feature_n = FeatureBuf_514;
         Mult_Buf[24].Weight_n = Wgt_9_514;
         Mult_Buf[25].Feature_n = FeatureBuf_515;
         Mult_Buf[25].Weight_n = Wgt_9_515;
         Mult_Buf[26].Feature_n = FeatureBuf_516;
         Mult_Buf[26].Weight_n = Wgt_9_516;
         Mult_Buf[27].Feature_n = FeatureBuf_517;
         Mult_Buf[27].Weight_n = Wgt_9_517;
         Mult_Buf[28].Feature_n = FeatureBuf_518;
         Mult_Buf[28].Weight_n = Wgt_9_518;
         Mult_Buf[29].Feature_n = FeatureBuf_519;
         Mult_Buf[29].Weight_n = Wgt_9_519;
         Mult_Buf[30].Feature_n = FeatureBuf_520;
         Mult_Buf[30].Weight_n = Wgt_9_520;
         Mult_Buf[31].Feature_n = FeatureBuf_521;
         Mult_Buf[31].Weight_n = Wgt_9_521;
         Mult_Buf[32].Feature_n = FeatureBuf_522;
         Mult_Buf[32].Weight_n = Wgt_9_522;
         Mult_Buf[33].Feature_n = FeatureBuf_523;
         Mult_Buf[33].Weight_n = Wgt_9_523;
         Mult_Buf[34].Feature_n = FeatureBuf_524;
         Mult_Buf[34].Weight_n = Wgt_9_524;
         Mult_Buf[35].Feature_n = FeatureBuf_525;
         Mult_Buf[35].Weight_n = Wgt_9_525;
         Mult_Buf[36].Feature_n = FeatureBuf_526;
         Mult_Buf[36].Weight_n = Wgt_9_526;
         Mult_Buf[37].Feature_n = FeatureBuf_527;
         Mult_Buf[37].Weight_n = Wgt_9_527;
         Mult_Buf[38].Feature_n = FeatureBuf_528;
         Mult_Buf[38].Weight_n = Wgt_9_528;
         Mult_Buf[39].Feature_n = FeatureBuf_529;
         Mult_Buf[39].Weight_n = Wgt_9_529;
         Mult_Buf[40].Feature_n = FeatureBuf_530;
         Mult_Buf[40].Weight_n = Wgt_9_530;
         Mult_Buf[41].Feature_n = FeatureBuf_531;
         Mult_Buf[41].Weight_n = Wgt_9_531;
         Mult_Buf[42].Feature_n = FeatureBuf_532;
         Mult_Buf[42].Weight_n = Wgt_9_532;
         Mult_Buf[43].Feature_n = FeatureBuf_533;
         Mult_Buf[43].Weight_n = Wgt_9_533;
         Mult_Buf[44].Feature_n = FeatureBuf_534;
         Mult_Buf[44].Weight_n = Wgt_9_534;
         Mult_Buf[45].Feature_n = FeatureBuf_535;
         Mult_Buf[45].Weight_n = Wgt_9_535;
         Mult_Buf[46].Feature_n = FeatureBuf_536;
         Mult_Buf[46].Weight_n = Wgt_9_536;
         Mult_Buf[47].Feature_n = FeatureBuf_537;
         Mult_Buf[47].Weight_n = Wgt_9_537;
         Mult_Buf[48].Feature_n = FeatureBuf_538;
         Mult_Buf[48].Weight_n = Wgt_9_538;
         Mult_Buf[49].Feature_n = FeatureBuf_539;
         Mult_Buf[49].Weight_n = Wgt_9_539;
         Mult_Buf[50].Feature_n = FeatureBuf_540;
         Mult_Buf[50].Weight_n = Wgt_9_540;
         Mult_Buf[51].Feature_n = FeatureBuf_541;
         Mult_Buf[51].Weight_n = Wgt_9_541;
         Mult_Buf[52].Feature_n = FeatureBuf_542;
         Mult_Buf[52].Weight_n = Wgt_9_542;
         Mult_Buf[53].Feature_n = FeatureBuf_543;
         Mult_Buf[53].Weight_n = Wgt_9_543;
         Mult_Buf[54].Feature_n = FeatureBuf_544;
         Mult_Buf[54].Weight_n = Wgt_9_544;
         Mult_Buf[55].Feature_n = FeatureBuf_545;
         Mult_Buf[55].Weight_n = Wgt_9_545;
         Mult_Buf[56].Feature_n = FeatureBuf_546;
         Mult_Buf[56].Weight_n = Wgt_9_546;
         Mult_Buf[57].Feature_n = FeatureBuf_547;
         Mult_Buf[57].Weight_n = Wgt_9_547;
         Mult_Buf[58].Feature_n = FeatureBuf_548;
         Mult_Buf[58].Weight_n = Wgt_9_548;
         Mult_Buf[59].Feature_n = FeatureBuf_549;
         Mult_Buf[59].Weight_n = Wgt_9_549;
         Mult_Buf[60].Feature_n = FeatureBuf_550;
         Mult_Buf[60].Weight_n = Wgt_9_550;
         Mult_Buf[61].Feature_n = FeatureBuf_551;
         Mult_Buf[61].Weight_n = Wgt_9_551;
         Mult_Buf[62].Feature_n = FeatureBuf_552;
         Mult_Buf[62].Weight_n = Wgt_9_552;
         Mult_Buf[63].Feature_n = FeatureBuf_553;
         Mult_Buf[63].Weight_n = Wgt_9_553;
         Mult_Buf[64].Feature_n = FeatureBuf_554;
         Mult_Buf[64].Weight_n = Wgt_9_554;
         Mult_Buf[65].Feature_n = FeatureBuf_555;
         Mult_Buf[65].Weight_n = Wgt_9_555;
         Mult_Buf[66].Feature_n = FeatureBuf_556;
         Mult_Buf[66].Weight_n = Wgt_9_556;
         Mult_Buf[67].Feature_n = FeatureBuf_557;
         Mult_Buf[67].Weight_n = Wgt_9_557;
         Mult_Buf[68].Feature_n = FeatureBuf_558;
         Mult_Buf[68].Weight_n = Wgt_9_558;
         Mult_Buf[69].Feature_n = FeatureBuf_559;
         Mult_Buf[69].Weight_n = Wgt_9_559;
         Mult_Buf[70].Feature_n = FeatureBuf_560;
         Mult_Buf[70].Weight_n = Wgt_9_560;
         Mult_Buf[71].Feature_n = FeatureBuf_561;
         Mult_Buf[71].Weight_n = Wgt_9_561;
         Mult_Buf[72].Feature_n = FeatureBuf_562;
         Mult_Buf[72].Weight_n = Wgt_9_562;
         Mult_Buf[73].Feature_n = FeatureBuf_563;
         Mult_Buf[73].Weight_n = Wgt_9_563;
         Mult_Buf[74].Feature_n = FeatureBuf_564;
         Mult_Buf[74].Weight_n = Wgt_9_564;
         Mult_Buf[75].Feature_n = FeatureBuf_565;
         Mult_Buf[75].Weight_n = Wgt_9_565;
         Mult_Buf[76].Feature_n = FeatureBuf_566;
         Mult_Buf[76].Weight_n = Wgt_9_566;
         Mult_Buf[77].Feature_n = FeatureBuf_567;
         Mult_Buf[77].Weight_n = Wgt_9_567;
         Mult_Buf[78].Feature_n = FeatureBuf_568;
         Mult_Buf[78].Weight_n = Wgt_9_568;
         Mult_Buf[79].Feature_n = FeatureBuf_569;
         Mult_Buf[79].Weight_n = Wgt_9_569;
         Mult_Buf[80].Feature_n = FeatureBuf_570;
         Mult_Buf[80].Weight_n = Wgt_9_570;
         Mult_Buf[81].Feature_n = FeatureBuf_571;
         Mult_Buf[81].Weight_n = Wgt_9_571;
         Mult_Buf[82].Feature_n = FeatureBuf_572;
         Mult_Buf[82].Weight_n = Wgt_9_572;
         Mult_Buf[83].Feature_n = FeatureBuf_573;
         Mult_Buf[83].Weight_n = Wgt_9_573;
         Mult_Buf[84].Feature_n = FeatureBuf_574;
         Mult_Buf[84].Weight_n = Wgt_9_574;
         Mult_Buf[85].Feature_n = FeatureBuf_575;
         Mult_Buf[85].Weight_n = Wgt_9_575;
         Mult_Buf[86].Feature_n = FeatureBuf_576;
         Mult_Buf[86].Weight_n = Wgt_9_576;
         Mult_Buf[87].Feature_n = FeatureBuf_577;
         Mult_Buf[87].Weight_n = Wgt_9_577;
         Mult_Buf[88].Feature_n = FeatureBuf_578;
         Mult_Buf[88].Weight_n = Wgt_9_578;
         Mult_Buf[89].Feature_n = FeatureBuf_579;
         Mult_Buf[89].Weight_n = Wgt_9_579;
         Mult_Buf[90].Feature_n = FeatureBuf_580;
         Mult_Buf[90].Weight_n = Wgt_9_580;
         Mult_Buf[91].Feature_n = FeatureBuf_581;
         Mult_Buf[91].Weight_n = Wgt_9_581;
         Mult_Buf[92].Feature_n = FeatureBuf_582;
         Mult_Buf[92].Weight_n = Wgt_9_582;
         Mult_Buf[93].Feature_n = FeatureBuf_583;
         Mult_Buf[93].Weight_n = Wgt_9_583;
         Mult_Buf[94].Feature_n = FeatureBuf_584;
         Mult_Buf[94].Weight_n = Wgt_9_584;
         Mult_Buf[95].Feature_n = FeatureBuf_585;
         Mult_Buf[95].Weight_n = Wgt_9_585;
         Mult_Buf[96].Feature_n = FeatureBuf_586;
         Mult_Buf[96].Weight_n = Wgt_9_586;
         Mult_Buf[97].Feature_n = FeatureBuf_587;
         Mult_Buf[97].Weight_n = Wgt_9_587;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     //Collect Partial result form Adder
         Res_6_7_n = Part_Res;
     //Feed to final Adder
         A1 = Part_Res;
         A2 = Res_6_6_n;
         A3 = Res_6_5_n;
         A4 = Res_6_4_n;
         A5 = Res_6_3_n;
         A6 = Res_6_2_n;
         A7 = Res_6_1_n;
         A8 = Res_6_0_n;
     end
    80:begin
     nxt_state = 81;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_588;
         Mult_Buf[0].Weight_n = Wgt_9_588;
         Mult_Buf[1].Feature_n = FeatureBuf_589;
         Mult_Buf[1].Weight_n = Wgt_9_589;
         Mult_Buf[2].Feature_n = FeatureBuf_590;
         Mult_Buf[2].Weight_n = Wgt_9_590;
         Mult_Buf[3].Feature_n = FeatureBuf_591;
         Mult_Buf[3].Weight_n = Wgt_9_591;
         Mult_Buf[4].Feature_n = FeatureBuf_592;
         Mult_Buf[4].Weight_n = Wgt_9_592;
         Mult_Buf[5].Feature_n = FeatureBuf_593;
         Mult_Buf[5].Weight_n = Wgt_9_593;
         Mult_Buf[6].Feature_n = FeatureBuf_594;
         Mult_Buf[6].Weight_n = Wgt_9_594;
         Mult_Buf[7].Feature_n = FeatureBuf_595;
         Mult_Buf[7].Weight_n = Wgt_9_595;
         Mult_Buf[8].Feature_n = FeatureBuf_596;
         Mult_Buf[8].Weight_n = Wgt_9_596;
         Mult_Buf[9].Feature_n = FeatureBuf_597;
         Mult_Buf[9].Weight_n = Wgt_9_597;
         Mult_Buf[10].Feature_n = FeatureBuf_598;
         Mult_Buf[10].Weight_n = Wgt_9_598;
         Mult_Buf[11].Feature_n = FeatureBuf_599;
         Mult_Buf[11].Weight_n = Wgt_9_599;
         Mult_Buf[12].Feature_n = FeatureBuf_600;
         Mult_Buf[12].Weight_n = Wgt_9_600;
         Mult_Buf[13].Feature_n = FeatureBuf_601;
         Mult_Buf[13].Weight_n = Wgt_9_601;
         Mult_Buf[14].Feature_n = FeatureBuf_602;
         Mult_Buf[14].Weight_n = Wgt_9_602;
         Mult_Buf[15].Feature_n = FeatureBuf_603;
         Mult_Buf[15].Weight_n = Wgt_9_603;
         Mult_Buf[16].Feature_n = FeatureBuf_604;
         Mult_Buf[16].Weight_n = Wgt_9_604;
         Mult_Buf[17].Feature_n = FeatureBuf_605;
         Mult_Buf[17].Weight_n = Wgt_9_605;
         Mult_Buf[18].Feature_n = FeatureBuf_606;
         Mult_Buf[18].Weight_n = Wgt_9_606;
         Mult_Buf[19].Feature_n = FeatureBuf_607;
         Mult_Buf[19].Weight_n = Wgt_9_607;
         Mult_Buf[20].Feature_n = FeatureBuf_608;
         Mult_Buf[20].Weight_n = Wgt_9_608;
         Mult_Buf[21].Feature_n = FeatureBuf_609;
         Mult_Buf[21].Weight_n = Wgt_9_609;
         Mult_Buf[22].Feature_n = FeatureBuf_610;
         Mult_Buf[22].Weight_n = Wgt_9_610;
         Mult_Buf[23].Feature_n = FeatureBuf_611;
         Mult_Buf[23].Weight_n = Wgt_9_611;
         Mult_Buf[24].Feature_n = FeatureBuf_612;
         Mult_Buf[24].Weight_n = Wgt_9_612;
         Mult_Buf[25].Feature_n = FeatureBuf_613;
         Mult_Buf[25].Weight_n = Wgt_9_613;
         Mult_Buf[26].Feature_n = FeatureBuf_614;
         Mult_Buf[26].Weight_n = Wgt_9_614;
         Mult_Buf[27].Feature_n = FeatureBuf_615;
         Mult_Buf[27].Weight_n = Wgt_9_615;
         Mult_Buf[28].Feature_n = FeatureBuf_616;
         Mult_Buf[28].Weight_n = Wgt_9_616;
         Mult_Buf[29].Feature_n = FeatureBuf_617;
         Mult_Buf[29].Weight_n = Wgt_9_617;
         Mult_Buf[30].Feature_n = FeatureBuf_618;
         Mult_Buf[30].Weight_n = Wgt_9_618;
         Mult_Buf[31].Feature_n = FeatureBuf_619;
         Mult_Buf[31].Weight_n = Wgt_9_619;
         Mult_Buf[32].Feature_n = FeatureBuf_620;
         Mult_Buf[32].Weight_n = Wgt_9_620;
         Mult_Buf[33].Feature_n = FeatureBuf_621;
         Mult_Buf[33].Weight_n = Wgt_9_621;
         Mult_Buf[34].Feature_n = FeatureBuf_622;
         Mult_Buf[34].Weight_n = Wgt_9_622;
         Mult_Buf[35].Feature_n = FeatureBuf_623;
         Mult_Buf[35].Weight_n = Wgt_9_623;
         Mult_Buf[36].Feature_n = FeatureBuf_624;
         Mult_Buf[36].Weight_n = Wgt_9_624;
         Mult_Buf[37].Feature_n = FeatureBuf_625;
         Mult_Buf[37].Weight_n = Wgt_9_625;
         Mult_Buf[38].Feature_n = FeatureBuf_626;
         Mult_Buf[38].Weight_n = Wgt_9_626;
         Mult_Buf[39].Feature_n = FeatureBuf_627;
         Mult_Buf[39].Weight_n = Wgt_9_627;
         Mult_Buf[40].Feature_n = FeatureBuf_628;
         Mult_Buf[40].Weight_n = Wgt_9_628;
         Mult_Buf[41].Feature_n = FeatureBuf_629;
         Mult_Buf[41].Weight_n = Wgt_9_629;
         Mult_Buf[42].Feature_n = FeatureBuf_630;
         Mult_Buf[42].Weight_n = Wgt_9_630;
         Mult_Buf[43].Feature_n = FeatureBuf_631;
         Mult_Buf[43].Weight_n = Wgt_9_631;
         Mult_Buf[44].Feature_n = FeatureBuf_632;
         Mult_Buf[44].Weight_n = Wgt_9_632;
         Mult_Buf[45].Feature_n = FeatureBuf_633;
         Mult_Buf[45].Weight_n = Wgt_9_633;
         Mult_Buf[46].Feature_n = FeatureBuf_634;
         Mult_Buf[46].Weight_n = Wgt_9_634;
         Mult_Buf[47].Feature_n = FeatureBuf_635;
         Mult_Buf[47].Weight_n = Wgt_9_635;
         Mult_Buf[48].Feature_n = FeatureBuf_636;
         Mult_Buf[48].Weight_n = Wgt_9_636;
         Mult_Buf[49].Feature_n = FeatureBuf_637;
         Mult_Buf[49].Weight_n = Wgt_9_637;
         Mult_Buf[50].Feature_n = FeatureBuf_638;
         Mult_Buf[50].Weight_n = Wgt_9_638;
         Mult_Buf[51].Feature_n = FeatureBuf_639;
         Mult_Buf[51].Weight_n = Wgt_9_639;
         Mult_Buf[52].Feature_n = FeatureBuf_640;
         Mult_Buf[52].Weight_n = Wgt_9_640;
         Mult_Buf[53].Feature_n = FeatureBuf_641;
         Mult_Buf[53].Weight_n = Wgt_9_641;
         Mult_Buf[54].Feature_n = FeatureBuf_642;
         Mult_Buf[54].Weight_n = Wgt_9_642;
         Mult_Buf[55].Feature_n = FeatureBuf_643;
         Mult_Buf[55].Weight_n = Wgt_9_643;
         Mult_Buf[56].Feature_n = FeatureBuf_644;
         Mult_Buf[56].Weight_n = Wgt_9_644;
         Mult_Buf[57].Feature_n = FeatureBuf_645;
         Mult_Buf[57].Weight_n = Wgt_9_645;
         Mult_Buf[58].Feature_n = FeatureBuf_646;
         Mult_Buf[58].Weight_n = Wgt_9_646;
         Mult_Buf[59].Feature_n = FeatureBuf_647;
         Mult_Buf[59].Weight_n = Wgt_9_647;
         Mult_Buf[60].Feature_n = FeatureBuf_648;
         Mult_Buf[60].Weight_n = Wgt_9_648;
         Mult_Buf[61].Feature_n = FeatureBuf_649;
         Mult_Buf[61].Weight_n = Wgt_9_649;
         Mult_Buf[62].Feature_n = FeatureBuf_650;
         Mult_Buf[62].Weight_n = Wgt_9_650;
         Mult_Buf[63].Feature_n = FeatureBuf_651;
         Mult_Buf[63].Weight_n = Wgt_9_651;
         Mult_Buf[64].Feature_n = FeatureBuf_652;
         Mult_Buf[64].Weight_n = Wgt_9_652;
         Mult_Buf[65].Feature_n = FeatureBuf_653;
         Mult_Buf[65].Weight_n = Wgt_9_653;
         Mult_Buf[66].Feature_n = FeatureBuf_654;
         Mult_Buf[66].Weight_n = Wgt_9_654;
         Mult_Buf[67].Feature_n = FeatureBuf_655;
         Mult_Buf[67].Weight_n = Wgt_9_655;
         Mult_Buf[68].Feature_n = FeatureBuf_656;
         Mult_Buf[68].Weight_n = Wgt_9_656;
         Mult_Buf[69].Feature_n = FeatureBuf_657;
         Mult_Buf[69].Weight_n = Wgt_9_657;
         Mult_Buf[70].Feature_n = FeatureBuf_658;
         Mult_Buf[70].Weight_n = Wgt_9_658;
         Mult_Buf[71].Feature_n = FeatureBuf_659;
         Mult_Buf[71].Weight_n = Wgt_9_659;
         Mult_Buf[72].Feature_n = FeatureBuf_660;
         Mult_Buf[72].Weight_n = Wgt_9_660;
         Mult_Buf[73].Feature_n = FeatureBuf_661;
         Mult_Buf[73].Weight_n = Wgt_9_661;
         Mult_Buf[74].Feature_n = FeatureBuf_662;
         Mult_Buf[74].Weight_n = Wgt_9_662;
         Mult_Buf[75].Feature_n = FeatureBuf_663;
         Mult_Buf[75].Weight_n = Wgt_9_663;
         Mult_Buf[76].Feature_n = FeatureBuf_664;
         Mult_Buf[76].Weight_n = Wgt_9_664;
         Mult_Buf[77].Feature_n = FeatureBuf_665;
         Mult_Buf[77].Weight_n = Wgt_9_665;
         Mult_Buf[78].Feature_n = FeatureBuf_666;
         Mult_Buf[78].Weight_n = Wgt_9_666;
         Mult_Buf[79].Feature_n = FeatureBuf_667;
         Mult_Buf[79].Weight_n = Wgt_9_667;
         Mult_Buf[80].Feature_n = FeatureBuf_668;
         Mult_Buf[80].Weight_n = Wgt_9_668;
         Mult_Buf[81].Feature_n = FeatureBuf_669;
         Mult_Buf[81].Weight_n = Wgt_9_669;
         Mult_Buf[82].Feature_n = FeatureBuf_670;
         Mult_Buf[82].Weight_n = Wgt_9_670;
         Mult_Buf[83].Feature_n = FeatureBuf_671;
         Mult_Buf[83].Weight_n = Wgt_9_671;
         Mult_Buf[84].Feature_n = FeatureBuf_672;
         Mult_Buf[84].Weight_n = Wgt_9_672;
         Mult_Buf[85].Feature_n = FeatureBuf_673;
         Mult_Buf[85].Weight_n = Wgt_9_673;
         Mult_Buf[86].Feature_n = FeatureBuf_674;
         Mult_Buf[86].Weight_n = Wgt_9_674;
         Mult_Buf[87].Feature_n = FeatureBuf_675;
         Mult_Buf[87].Weight_n = Wgt_9_675;
         Mult_Buf[88].Feature_n = FeatureBuf_676;
         Mult_Buf[88].Weight_n = Wgt_9_676;
         Mult_Buf[89].Feature_n = FeatureBuf_677;
         Mult_Buf[89].Weight_n = Wgt_9_677;
         Mult_Buf[90].Feature_n = FeatureBuf_678;
         Mult_Buf[90].Weight_n = Wgt_9_678;
         Mult_Buf[91].Feature_n = FeatureBuf_679;
         Mult_Buf[91].Weight_n = Wgt_9_679;
         Mult_Buf[92].Feature_n = FeatureBuf_680;
         Mult_Buf[92].Weight_n = Wgt_9_680;
         Mult_Buf[93].Feature_n = FeatureBuf_681;
         Mult_Buf[93].Weight_n = Wgt_9_681;
         Mult_Buf[94].Feature_n = FeatureBuf_682;
         Mult_Buf[94].Weight_n = Wgt_9_682;
         Mult_Buf[95].Feature_n = FeatureBuf_683;
         Mult_Buf[95].Weight_n = Wgt_9_683;
         Mult_Buf[96].Feature_n = FeatureBuf_684;
         Mult_Buf[96].Weight_n = Wgt_9_684;
         Mult_Buf[97].Feature_n = FeatureBuf_685;
         Mult_Buf[97].Weight_n = Wgt_9_685;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     //Collect Partial result form Adder
         Res_7_0_n = Part_Res;
     end
    81:begin
     nxt_state = 82;
     //Feed input to Multipliers
         Mult_Buf[0].Feature_n = FeatureBuf_686;
         Mult_Buf[0].Weight_n = Wgt_9_686;
         Mult_Buf[1].Feature_n = FeatureBuf_687;
         Mult_Buf[1].Weight_n = Wgt_9_687;
         Mult_Buf[2].Feature_n = FeatureBuf_688;
         Mult_Buf[2].Weight_n = Wgt_9_688;
         Mult_Buf[3].Feature_n = FeatureBuf_689;
         Mult_Buf[3].Weight_n = Wgt_9_689;
         Mult_Buf[4].Feature_n = FeatureBuf_690;
         Mult_Buf[4].Weight_n = Wgt_9_690;
         Mult_Buf[5].Feature_n = FeatureBuf_691;
         Mult_Buf[5].Weight_n = Wgt_9_691;
         Mult_Buf[6].Feature_n = FeatureBuf_692;
         Mult_Buf[6].Weight_n = Wgt_9_692;
         Mult_Buf[7].Feature_n = FeatureBuf_693;
         Mult_Buf[7].Weight_n = Wgt_9_693;
         Mult_Buf[8].Feature_n = FeatureBuf_694;
         Mult_Buf[8].Weight_n = Wgt_9_694;
         Mult_Buf[9].Feature_n = FeatureBuf_695;
         Mult_Buf[9].Weight_n = Wgt_9_695;
         Mult_Buf[10].Feature_n = FeatureBuf_696;
         Mult_Buf[10].Weight_n = Wgt_9_696;
         Mult_Buf[11].Feature_n = FeatureBuf_697;
         Mult_Buf[11].Weight_n = Wgt_9_697;
         Mult_Buf[12].Feature_n = FeatureBuf_698;
         Mult_Buf[12].Weight_n = Wgt_9_698;
         Mult_Buf[13].Feature_n = FeatureBuf_699;
         Mult_Buf[13].Weight_n = Wgt_9_699;
         Mult_Buf[14].Feature_n = FeatureBuf_700;
         Mult_Buf[14].Weight_n = Wgt_9_700;
         Mult_Buf[15].Feature_n = FeatureBuf_701;
         Mult_Buf[15].Weight_n = Wgt_9_701;
         Mult_Buf[16].Feature_n = FeatureBuf_702;
         Mult_Buf[16].Weight_n = Wgt_9_702;
         Mult_Buf[17].Feature_n = FeatureBuf_703;
         Mult_Buf[17].Weight_n = Wgt_9_703;
         Mult_Buf[18].Feature_n = FeatureBuf_704;
         Mult_Buf[18].Weight_n = Wgt_9_704;
         Mult_Buf[19].Feature_n = FeatureBuf_705;
         Mult_Buf[19].Weight_n = Wgt_9_705;
         Mult_Buf[20].Feature_n = FeatureBuf_706;
         Mult_Buf[20].Weight_n = Wgt_9_706;
         Mult_Buf[21].Feature_n = FeatureBuf_707;
         Mult_Buf[21].Weight_n = Wgt_9_707;
         Mult_Buf[22].Feature_n = FeatureBuf_708;
         Mult_Buf[22].Weight_n = Wgt_9_708;
         Mult_Buf[23].Feature_n = FeatureBuf_709;
         Mult_Buf[23].Weight_n = Wgt_9_709;
         Mult_Buf[24].Feature_n = FeatureBuf_710;
         Mult_Buf[24].Weight_n = Wgt_9_710;
         Mult_Buf[25].Feature_n = FeatureBuf_711;
         Mult_Buf[25].Weight_n = Wgt_9_711;
         Mult_Buf[26].Feature_n = FeatureBuf_712;
         Mult_Buf[26].Weight_n = Wgt_9_712;
         Mult_Buf[27].Feature_n = FeatureBuf_713;
         Mult_Buf[27].Weight_n = Wgt_9_713;
         Mult_Buf[28].Feature_n = FeatureBuf_714;
         Mult_Buf[28].Weight_n = Wgt_9_714;
         Mult_Buf[29].Feature_n = FeatureBuf_715;
         Mult_Buf[29].Weight_n = Wgt_9_715;
         Mult_Buf[30].Feature_n = FeatureBuf_716;
         Mult_Buf[30].Weight_n = Wgt_9_716;
         Mult_Buf[31].Feature_n = FeatureBuf_717;
         Mult_Buf[31].Weight_n = Wgt_9_717;
         Mult_Buf[32].Feature_n = FeatureBuf_718;
         Mult_Buf[32].Weight_n = Wgt_9_718;
         Mult_Buf[33].Feature_n = FeatureBuf_719;
         Mult_Buf[33].Weight_n = Wgt_9_719;
         Mult_Buf[34].Feature_n = FeatureBuf_720;
         Mult_Buf[34].Weight_n = Wgt_9_720;
         Mult_Buf[35].Feature_n = FeatureBuf_721;
         Mult_Buf[35].Weight_n = Wgt_9_721;
         Mult_Buf[36].Feature_n = FeatureBuf_722;
         Mult_Buf[36].Weight_n = Wgt_9_722;
         Mult_Buf[37].Feature_n = FeatureBuf_723;
         Mult_Buf[37].Weight_n = Wgt_9_723;
         Mult_Buf[38].Feature_n = FeatureBuf_724;
         Mult_Buf[38].Weight_n = Wgt_9_724;
         Mult_Buf[39].Feature_n = FeatureBuf_725;
         Mult_Buf[39].Weight_n = Wgt_9_725;
         Mult_Buf[40].Feature_n = FeatureBuf_726;
         Mult_Buf[40].Weight_n = Wgt_9_726;
         Mult_Buf[41].Feature_n = FeatureBuf_727;
         Mult_Buf[41].Weight_n = Wgt_9_727;
         Mult_Buf[42].Feature_n = FeatureBuf_728;
         Mult_Buf[42].Weight_n = Wgt_9_728;
         Mult_Buf[43].Feature_n = FeatureBuf_729;
         Mult_Buf[43].Weight_n = Wgt_9_729;
         Mult_Buf[44].Feature_n = FeatureBuf_730;
         Mult_Buf[44].Weight_n = Wgt_9_730;
         Mult_Buf[45].Feature_n = FeatureBuf_731;
         Mult_Buf[45].Weight_n = Wgt_9_731;
         Mult_Buf[46].Feature_n = FeatureBuf_732;
         Mult_Buf[46].Weight_n = Wgt_9_732;
         Mult_Buf[47].Feature_n = FeatureBuf_733;
         Mult_Buf[47].Weight_n = Wgt_9_733;
         Mult_Buf[48].Feature_n = FeatureBuf_734;
         Mult_Buf[48].Weight_n = Wgt_9_734;
         Mult_Buf[49].Feature_n = FeatureBuf_735;
         Mult_Buf[49].Weight_n = Wgt_9_735;
         Mult_Buf[50].Feature_n = FeatureBuf_736;
         Mult_Buf[50].Weight_n = Wgt_9_736;
         Mult_Buf[51].Feature_n = FeatureBuf_737;
         Mult_Buf[51].Weight_n = Wgt_9_737;
         Mult_Buf[52].Feature_n = FeatureBuf_738;
         Mult_Buf[52].Weight_n = Wgt_9_738;
         Mult_Buf[53].Feature_n = FeatureBuf_739;
         Mult_Buf[53].Weight_n = Wgt_9_739;
         Mult_Buf[54].Feature_n = FeatureBuf_740;
         Mult_Buf[54].Weight_n = Wgt_9_740;
         Mult_Buf[55].Feature_n = FeatureBuf_741;
         Mult_Buf[55].Weight_n = Wgt_9_741;
         Mult_Buf[56].Feature_n = FeatureBuf_742;
         Mult_Buf[56].Weight_n = Wgt_9_742;
         Mult_Buf[57].Feature_n = FeatureBuf_743;
         Mult_Buf[57].Weight_n = Wgt_9_743;
         Mult_Buf[58].Feature_n = FeatureBuf_744;
         Mult_Buf[58].Weight_n = Wgt_9_744;
         Mult_Buf[59].Feature_n = FeatureBuf_745;
         Mult_Buf[59].Weight_n = Wgt_9_745;
         Mult_Buf[60].Feature_n = FeatureBuf_746;
         Mult_Buf[60].Weight_n = Wgt_9_746;
         Mult_Buf[61].Feature_n = FeatureBuf_747;
         Mult_Buf[61].Weight_n = Wgt_9_747;
         Mult_Buf[62].Feature_n = FeatureBuf_748;
         Mult_Buf[62].Weight_n = Wgt_9_748;
         Mult_Buf[63].Feature_n = FeatureBuf_749;
         Mult_Buf[63].Weight_n = Wgt_9_749;
         Mult_Buf[64].Feature_n = FeatureBuf_750;
         Mult_Buf[64].Weight_n = Wgt_9_750;
         Mult_Buf[65].Feature_n = FeatureBuf_751;
         Mult_Buf[65].Weight_n = Wgt_9_751;
         Mult_Buf[66].Feature_n = FeatureBuf_752;
         Mult_Buf[66].Weight_n = Wgt_9_752;
         Mult_Buf[67].Feature_n = FeatureBuf_753;
         Mult_Buf[67].Weight_n = Wgt_9_753;
         Mult_Buf[68].Feature_n = FeatureBuf_754;
         Mult_Buf[68].Weight_n = Wgt_9_754;
         Mult_Buf[69].Feature_n = FeatureBuf_755;
         Mult_Buf[69].Weight_n = Wgt_9_755;
         Mult_Buf[70].Feature_n = FeatureBuf_756;
         Mult_Buf[70].Weight_n = Wgt_9_756;
         Mult_Buf[71].Feature_n = FeatureBuf_757;
         Mult_Buf[71].Weight_n = Wgt_9_757;
         Mult_Buf[72].Feature_n = FeatureBuf_758;
         Mult_Buf[72].Weight_n = Wgt_9_758;
         Mult_Buf[73].Feature_n = FeatureBuf_759;
         Mult_Buf[73].Weight_n = Wgt_9_759;
         Mult_Buf[74].Feature_n = FeatureBuf_760;
         Mult_Buf[74].Weight_n = Wgt_9_760;
         Mult_Buf[75].Feature_n = FeatureBuf_761;
         Mult_Buf[75].Weight_n = Wgt_9_761;
         Mult_Buf[76].Feature_n = FeatureBuf_762;
         Mult_Buf[76].Weight_n = Wgt_9_762;
         Mult_Buf[77].Feature_n = FeatureBuf_763;
         Mult_Buf[77].Weight_n = Wgt_9_763;
         Mult_Buf[78].Feature_n = FeatureBuf_764;
         Mult_Buf[78].Weight_n = Wgt_9_764;
         Mult_Buf[79].Feature_n = FeatureBuf_765;
         Mult_Buf[79].Weight_n = Wgt_9_765;
         Mult_Buf[80].Feature_n = FeatureBuf_766;
         Mult_Buf[80].Weight_n = Wgt_9_766;
         Mult_Buf[81].Feature_n = FeatureBuf_767;
         Mult_Buf[81].Weight_n = Wgt_9_767;
         Mult_Buf[82].Feature_n = FeatureBuf_768;
         Mult_Buf[82].Weight_n = Wgt_9_768;
         Mult_Buf[83].Feature_n = FeatureBuf_769;
         Mult_Buf[83].Weight_n = Wgt_9_769;
         Mult_Buf[84].Feature_n = FeatureBuf_770;
         Mult_Buf[84].Weight_n = Wgt_9_770;
         Mult_Buf[85].Feature_n = FeatureBuf_771;
         Mult_Buf[85].Weight_n = Wgt_9_771;
         Mult_Buf[86].Feature_n = FeatureBuf_772;
         Mult_Buf[86].Weight_n = Wgt_9_772;
         Mult_Buf[87].Feature_n = FeatureBuf_773;
         Mult_Buf[87].Weight_n = Wgt_9_773;
         Mult_Buf[88].Feature_n = FeatureBuf_774;
         Mult_Buf[88].Weight_n = Wgt_9_774;
         Mult_Buf[89].Feature_n = FeatureBuf_775;
         Mult_Buf[89].Weight_n = Wgt_9_775;
         Mult_Buf[90].Feature_n = FeatureBuf_776;
         Mult_Buf[90].Weight_n = Wgt_9_776;
         Mult_Buf[91].Feature_n = FeatureBuf_777;
         Mult_Buf[91].Weight_n = Wgt_9_777;
         Mult_Buf[92].Feature_n = FeatureBuf_778;
         Mult_Buf[92].Weight_n = Wgt_9_778;
         Mult_Buf[93].Feature_n = FeatureBuf_779;
         Mult_Buf[93].Weight_n = Wgt_9_779;
         Mult_Buf[94].Feature_n = FeatureBuf_780;
         Mult_Buf[94].Weight_n = Wgt_9_780;
         Mult_Buf[95].Feature_n = FeatureBuf_781;
         Mult_Buf[95].Weight_n = Wgt_9_781;
         Mult_Buf[96].Feature_n = FeatureBuf_782;
         Mult_Buf[96].Weight_n = Wgt_9_782;
         Mult_Buf[97].Feature_n = FeatureBuf_783;
         Mult_Buf[97].Weight_n = Wgt_9_783;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     //Collect Partial result form Adder
         Res_7_1_n = Part_Res;
     end
    82:begin
     nxt_state = 83;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     //Collect Partial result form Adder
         Res_7_2_n = Part_Res;
     end
    83:begin
     nxt_state = 84;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     //Collect Partial result form Adder
         Res_7_3_n = Part_Res;
     end
    84:begin
     nxt_state = 85;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     //Collect Partial result form Adder
         Res_7_4_n = Part_Res;
     end
    85:begin
     nxt_state = 86;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     //Collect Partial result form Adder
         Res_7_5_n = Part_Res;
     //Collect result from final Adder
         Res6_n = Final_Res;
     end
    86:begin
     nxt_state = 87;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     //Collect Partial result form Adder
         Res_7_6_n = Part_Res;
     end
    87:begin
     nxt_state = 88;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     //Collect Partial result form Adder
         Res_7_7_n = Part_Res;
     //Feed to final Adder
         A1 = Part_Res;
         A2 = Res_7_6_n;
         A3 = Res_7_5_n;
         A4 = Res_7_4_n;
         A5 = Res_7_3_n;
         A6 = Res_7_2_n;
         A7 = Res_7_1_n;
         A8 = Res_7_0_n;
     end
    88:begin
     nxt_state = 89;
     //Feed input to Adders
         Add_Buf[0].A_n = Multiplyer_matrix[0].Result;
         Add_Buf[0].B_n = Multiplyer_matrix[1].Result;
         Add_Buf[1].A_n = Multiplyer_matrix[2].Result;
         Add_Buf[1].B_n = Multiplyer_matrix[3].Result;
         Add_Buf[2].A_n = Multiplyer_matrix[4].Result;
         Add_Buf[2].B_n = Multiplyer_matrix[5].Result;
         Add_Buf[3].A_n = Multiplyer_matrix[6].Result;
         Add_Buf[3].B_n = Multiplyer_matrix[7].Result;
         Add_Buf[4].A_n = Multiplyer_matrix[8].Result;
         Add_Buf[4].B_n = Multiplyer_matrix[9].Result;
         Add_Buf[5].A_n = Multiplyer_matrix[10].Result;
         Add_Buf[5].B_n = Multiplyer_matrix[11].Result;
         Add_Buf[6].A_n = Multiplyer_matrix[12].Result;
         Add_Buf[6].B_n = Multiplyer_matrix[13].Result;
         Add_Buf[7].A_n = Multiplyer_matrix[14].Result;
         Add_Buf[7].B_n = Multiplyer_matrix[15].Result;
         Add_Buf[8].A_n = Multiplyer_matrix[16].Result;
         Add_Buf[8].B_n = Multiplyer_matrix[17].Result;
         Add_Buf[9].A_n = Multiplyer_matrix[18].Result;
         Add_Buf[9].B_n = Multiplyer_matrix[19].Result;
         Add_Buf[10].A_n = Multiplyer_matrix[20].Result;
         Add_Buf[10].B_n = Multiplyer_matrix[21].Result;
         Add_Buf[11].A_n = Multiplyer_matrix[22].Result;
         Add_Buf[11].B_n = Multiplyer_matrix[23].Result;
         Add_Buf[12].A_n = Multiplyer_matrix[24].Result;
         Add_Buf[12].B_n = Multiplyer_matrix[25].Result;
         Add_Buf[13].A_n = Multiplyer_matrix[26].Result;
         Add_Buf[13].B_n = Multiplyer_matrix[27].Result;
         Add_Buf[14].A_n = Multiplyer_matrix[28].Result;
         Add_Buf[14].B_n = Multiplyer_matrix[29].Result;
         Add_Buf[15].A_n = Multiplyer_matrix[30].Result;
         Add_Buf[15].B_n = Multiplyer_matrix[31].Result;
         Add_Buf[16].A_n = Multiplyer_matrix[32].Result;
         Add_Buf[16].B_n = Multiplyer_matrix[33].Result;
         Add_Buf[17].A_n = Multiplyer_matrix[34].Result;
         Add_Buf[17].B_n = Multiplyer_matrix[35].Result;
         Add_Buf[18].A_n = Multiplyer_matrix[36].Result;
         Add_Buf[18].B_n = Multiplyer_matrix[37].Result;
         Add_Buf[19].A_n = Multiplyer_matrix[38].Result;
         Add_Buf[19].B_n = Multiplyer_matrix[39].Result;
         Add_Buf[20].A_n = Multiplyer_matrix[40].Result;
         Add_Buf[20].B_n = Multiplyer_matrix[41].Result;
         Add_Buf[21].A_n = Multiplyer_matrix[42].Result;
         Add_Buf[21].B_n = Multiplyer_matrix[43].Result;
         Add_Buf[22].A_n = Multiplyer_matrix[44].Result;
         Add_Buf[22].B_n = Multiplyer_matrix[45].Result;
         Add_Buf[23].A_n = Multiplyer_matrix[46].Result;
         Add_Buf[23].B_n = Multiplyer_matrix[47].Result;
         Add_Buf[24].A_n = Multiplyer_matrix[48].Result;
         Add_Buf[24].B_n = Multiplyer_matrix[49].Result;
         Add_Buf[25].A_n = Multiplyer_matrix[50].Result;
         Add_Buf[25].B_n = Multiplyer_matrix[51].Result;
         Add_Buf[26].A_n = Multiplyer_matrix[52].Result;
         Add_Buf[26].B_n = Multiplyer_matrix[53].Result;
         Add_Buf[27].A_n = Multiplyer_matrix[54].Result;
         Add_Buf[27].B_n = Multiplyer_matrix[55].Result;
         Add_Buf[28].A_n = Multiplyer_matrix[56].Result;
         Add_Buf[28].B_n = Multiplyer_matrix[57].Result;
         Add_Buf[29].A_n = Multiplyer_matrix[58].Result;
         Add_Buf[29].B_n = Multiplyer_matrix[59].Result;
         Add_Buf[30].A_n = Multiplyer_matrix[60].Result;
         Add_Buf[30].B_n = Multiplyer_matrix[61].Result;
         Add_Buf[31].A_n = Multiplyer_matrix[62].Result;
         Add_Buf[31].B_n = Multiplyer_matrix[63].Result;
         Add_Buf[32].A_n = Multiplyer_matrix[64].Result;
         Add_Buf[32].B_n = Multiplyer_matrix[65].Result;
         Add_Buf[33].A_n = Multiplyer_matrix[66].Result;
         Add_Buf[33].B_n = Multiplyer_matrix[67].Result;
         Add_Buf[34].A_n = Multiplyer_matrix[68].Result;
         Add_Buf[34].B_n = Multiplyer_matrix[69].Result;
         Add_Buf[35].A_n = Multiplyer_matrix[70].Result;
         Add_Buf[35].B_n = Multiplyer_matrix[71].Result;
         Add_Buf[36].A_n = Multiplyer_matrix[72].Result;
         Add_Buf[36].B_n = Multiplyer_matrix[73].Result;
         Add_Buf[37].A_n = Multiplyer_matrix[74].Result;
         Add_Buf[37].B_n = Multiplyer_matrix[75].Result;
         Add_Buf[38].A_n = Multiplyer_matrix[76].Result;
         Add_Buf[38].B_n = Multiplyer_matrix[77].Result;
         Add_Buf[39].A_n = Multiplyer_matrix[78].Result;
         Add_Buf[39].B_n = Multiplyer_matrix[79].Result;
         Add_Buf[40].A_n = Multiplyer_matrix[80].Result;
         Add_Buf[40].B_n = Multiplyer_matrix[81].Result;
         Add_Buf[41].A_n = Multiplyer_matrix[82].Result;
         Add_Buf[41].B_n = Multiplyer_matrix[83].Result;
         Add_Buf[42].A_n = Multiplyer_matrix[84].Result;
         Add_Buf[42].B_n = Multiplyer_matrix[85].Result;
         Add_Buf[43].A_n = Multiplyer_matrix[86].Result;
         Add_Buf[43].B_n = Multiplyer_matrix[87].Result;
         Add_Buf[44].A_n = Multiplyer_matrix[88].Result;
         Add_Buf[44].B_n = Multiplyer_matrix[89].Result;
         Add_Buf[45].A_n = Multiplyer_matrix[90].Result;
         Add_Buf[45].B_n = Multiplyer_matrix[91].Result;
         Add_Buf[46].A_n = Multiplyer_matrix[92].Result;
         Add_Buf[46].B_n = Multiplyer_matrix[93].Result;
         Add_Buf[47].A_n = Multiplyer_matrix[94].Result;
         Add_Buf[47].B_n = Multiplyer_matrix[95].Result;
         Add_Buf[48].A_n = Multiplyer_matrix[96].Result;
         Add_Buf[48].B_n = Multiplyer_matrix[97].Result;
     //Collect Partial result form Adder
         Res_8_0_n = Part_Res;
     end
    89:begin
     nxt_state = 90;
     //Collect Partial result form Adder
         Res_8_1_n = Part_Res;
     end
    90:begin
     nxt_state = 91;
     //Collect Partial result form Adder
         Res_8_2_n = Part_Res;
     end
    91:begin
     nxt_state = 92;
     //Collect Partial result form Adder
         Res_8_3_n = Part_Res;
     end
    92:begin
     nxt_state = 93;
     //Collect Partial result form Adder
         Res_8_4_n = Part_Res;
     end
    93:begin
     nxt_state = 94;
     //Collect Partial result form Adder
         Res_8_5_n = Part_Res;
     //Collect result from final Adder
         Res7_n = Final_Res;
     end
    94:begin
     nxt_state = 95;
     //Collect Partial result form Adder
         Res_8_6_n = Part_Res;
     end
    95:begin
     nxt_state = 96;
     //Collect Partial result form Adder
         Res_8_7_n = Part_Res;
     //Feed to final Adder
         A1 = Part_Res;
         A2 = Res_8_6_n;
         A3 = Res_8_5_n;
         A4 = Res_8_4_n;
         A5 = Res_8_3_n;
         A6 = Res_8_2_n;
         A7 = Res_8_1_n;
         A8 = Res_8_0_n;
     end
    96:begin
     nxt_state = 97;
     //Collect Partial result form Adder
         Res_9_0_n = Part_Res;
     end
    97:begin
     nxt_state = 98;
     //Collect Partial result form Adder
         Res_9_1_n = Part_Res;
     end
    98:begin
     nxt_state = 99;
     //Collect Partial result form Adder
         Res_9_2_n = Part_Res;
     end
    99:begin
     nxt_state = 100;
     //Collect Partial result form Adder
         Res_9_3_n = Part_Res;
     end
    100:begin
     nxt_state = 101;
     //Collect Partial result form Adder
         Res_9_4_n = Part_Res;
     end
    101:begin
     nxt_state = 102;
     //Collect Partial result form Adder
         Res_9_5_n = Part_Res;
     //Collect result from final Adder
         Res8_n = Final_Res;
     end
    102:begin
     nxt_state = 103;
     //Collect Partial result form Adder
         Res_9_6_n = Part_Res;
     end
    103:begin
     nxt_state = 104;
     //Collect Partial result form Adder
         Res_9_7_n = Part_Res;
     //Feed to final Adder
         A1 = Part_Res;
         A2 = Res_9_6_n;
         A3 = Res_9_5_n;
         A4 = Res_9_4_n;
         A5 = Res_9_3_n;
         A6 = Res_9_2_n;
         A7 = Res_9_1_n;
         A8 = Res_9_0_n;
     end
    104:begin
     nxt_state = 105;
     end
    105:begin
     nxt_state = 106;
     end
    106:begin
     nxt_state = 107;
     end
    107:begin
     nxt_state = 108;
     end
    108:begin
     nxt_state = 109;
     end
    109:begin
     nxt_state = 110;
     //Collect result from final Adder
         Res9_n = Final_Res;
     end


///////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////
    110:begin
        // Add bias to the result
        Add_Buf[0].A_n = Res0;
        Add_Buf[0].B_n = {{7{Wgt_0_784[18]}},Wgt_0_784};
        Add_Buf[1].A_n = Res1;
        Add_Buf[1].B_n = {{7{Wgt_1_784[18]}},Wgt_1_784};
        Add_Buf[2].A_n = Res2;
        Add_Buf[2].B_n = {{7{Wgt_2_784[18]}},Wgt_2_784};
        Add_Buf[3].A_n = Res3;
        Add_Buf[3].B_n = {{7{Wgt_3_784[18]}},Wgt_3_784};
        Add_Buf[4].A_n = Res4;
        Add_Buf[4].B_n = {{7{Wgt_4_784[18]}},Wgt_4_784};
        Add_Buf[5].A_n = Res5;
        Add_Buf[5].B_n = {{7{Wgt_5_784[18]}},Wgt_5_784};
        Add_Buf[6].A_n = Res6;
        Add_Buf[6].B_n = {{7{Wgt_6_784[18]}},Wgt_6_784};
        Add_Buf[7].A_n = Res7;
        Add_Buf[7].B_n = {{7{Wgt_7_784[18]}},Wgt_7_784};
        Add_Buf[8].A_n = Res8;
        Add_Buf[8].B_n = {{7{Wgt_8_784[18]}},Wgt_8_784};
        Add_Buf[9].A_n = Res9;
        Add_Buf[9].B_n = {{7{Wgt_9_784[18]}},Wgt_9_784};
        nxt_state = 111;
    end

    111:begin
        // Wait for the bias calculation finish
        nxt_state = 112;
    end

    112: begin
        nxt_state = 113;
    end
    113:begin
        // Read final number
            Res0_n = Adder_Base[0].Res;
            Res1_n = Adder_Base[1].Res;
            Res2_n = Adder_Base[2].Res;
            Res3_n = Adder_Base[3].Res;
            Res4_n = Adder_Base[4].Res;
            Res5_n = Adder_Base[5].Res;
            Res6_n = Adder_Base[6].Res;
            Res7_n = Adder_Base[7].Res;
            Res8_n = Adder_Base[8].Res;
            Res9_n = Adder_Base[9].Res;
            nxt_state = 114;
    end

    114:begin
        // Start comparasion
        W11_n = Res0>Res1?0:1;
        W12_n = Res2>Res3?2:3;
        W13_n = Res4>Res5?4:5;
        W14_n = Res6>Res7?6:7;
        W15_n = Res8>Res9?8:9;
        V11_n = Res0>Res1?Res0:Res1;
        V12_n = Res2>Res3?Res2:Res3;
        V13_n = Res4>Res5?Res4:Res5;
        V14_n = Res6>Res7?Res6:Res7;
        V15_n = Res8>Res9?Res8:Res9;
        nxt_state = 115;
    end
    115:begin
        V15_n = V15;
        W15_n = W15;
        W21_n = V11>V12?W11:W12;
        W22_n = V13>V14?W13:W14;
        V21_n = V11>V12?V11:V12;
        V22_n = V13>V14?V13:V14;
        nxt_state = 116;
    end
    116:begin
        W31_n = V21>V22?W21:W22;
        W32_n = V21>V15?W21:W15;
        V31_n = V21>V22?V21:V22;
        V32_n = V21>V15?V21:V15;
        nxt_state = 117;
    end
    117:begin
        Output_Valid = 1;
        nxt_state =Input_Valid?1:118;
    end
    endcase
end
endmodule